magic
tech sky130A
magscale 1 2
timestamp 1693968996
<< viali >>
rect 1501 39049 1535 39083
rect 4905 39049 4939 39083
rect 9321 39049 9355 39083
rect 11621 39049 11655 39083
rect 13185 39049 13219 39083
rect 17785 39049 17819 39083
rect 22109 39049 22143 39083
rect 27169 39049 27203 39083
rect 33149 39049 33183 39083
rect 35725 39049 35759 39083
rect 11897 38981 11931 39015
rect 15761 38981 15795 39015
rect 31217 38981 31251 39015
rect 1777 38913 1811 38947
rect 5089 38913 5123 38947
rect 9229 38913 9263 38947
rect 12081 38913 12115 38947
rect 13001 38913 13035 38947
rect 17969 38913 18003 38947
rect 19441 38913 19475 38947
rect 20085 38913 20119 38947
rect 22385 38913 22419 38947
rect 27077 38913 27111 38947
rect 27721 38913 27755 38947
rect 33057 38913 33091 38947
rect 35633 38913 35667 38947
rect 37473 38913 37507 38947
rect 20361 38845 20395 38879
rect 15577 38777 15611 38811
rect 31033 38777 31067 38811
rect 37657 38777 37691 38811
rect 12265 38709 12299 38743
rect 19625 38709 19659 38743
rect 27629 38709 27663 38743
rect 4997 38505 5031 38539
rect 8769 38505 8803 38539
rect 18337 38505 18371 38539
rect 32229 38505 32263 38539
rect 34897 38505 34931 38539
rect 37841 38505 37875 38539
rect 11069 38369 11103 38403
rect 19533 38369 19567 38403
rect 27261 38369 27295 38403
rect 5181 38301 5215 38335
rect 8585 38301 8619 38335
rect 9045 38301 9079 38335
rect 9137 38301 9171 38335
rect 9321 38301 9355 38335
rect 13093 38301 13127 38335
rect 13277 38301 13311 38335
rect 13369 38301 13403 38335
rect 18521 38301 18555 38335
rect 18889 38301 18923 38335
rect 18981 38301 19015 38335
rect 19257 38301 19291 38335
rect 21281 38301 21315 38335
rect 21557 38301 21591 38335
rect 21649 38301 21683 38335
rect 21833 38301 21867 38335
rect 25053 38301 25087 38335
rect 25145 38301 25179 38335
rect 25329 38301 25363 38335
rect 29561 38301 29595 38335
rect 29653 38301 29687 38335
rect 32045 38301 32079 38335
rect 34713 38301 34747 38335
rect 9597 38233 9631 38267
rect 12817 38233 12851 38267
rect 22109 38233 22143 38267
rect 25605 38233 25639 38267
rect 27537 38233 27571 38267
rect 29285 38233 29319 38267
rect 37565 38233 37599 38267
rect 11345 38165 11379 38199
rect 21005 38165 21039 38199
rect 21465 38165 21499 38199
rect 23581 38165 23615 38199
rect 27077 38165 27111 38199
rect 9781 37961 9815 37995
rect 10241 37961 10275 37995
rect 12265 37961 12299 37995
rect 12357 37961 12391 37995
rect 19441 37961 19475 37995
rect 19809 37961 19843 37995
rect 22017 37961 22051 37995
rect 22477 37961 22511 37995
rect 24869 37961 24903 37995
rect 26249 37961 26283 37995
rect 26801 37961 26835 37995
rect 27905 37961 27939 37995
rect 10701 37893 10735 37927
rect 11805 37893 11839 37927
rect 11897 37893 11931 37927
rect 14039 37893 14073 37927
rect 14473 37893 14507 37927
rect 16681 37893 16715 37927
rect 17049 37893 17083 37927
rect 17417 37893 17451 37927
rect 23581 37893 23615 37927
rect 24409 37893 24443 37927
rect 25789 37893 25823 37927
rect 9965 37825 9999 37859
rect 10609 37825 10643 37859
rect 12541 37825 12575 37859
rect 13277 37825 13311 37859
rect 13737 37825 13771 37859
rect 13829 37825 13863 37859
rect 13921 37825 13955 37859
rect 14376 37825 14410 37859
rect 14565 37825 14599 37859
rect 14749 37825 14783 37859
rect 15945 37825 15979 37859
rect 16129 37825 16163 37859
rect 16221 37825 16255 37859
rect 16313 37825 16347 37859
rect 16865 37825 16899 37859
rect 17233 37825 17267 37859
rect 17509 37825 17543 37859
rect 17601 37825 17635 37859
rect 20361 37825 20395 37859
rect 20729 37825 20763 37859
rect 22385 37825 22419 37859
rect 23397 37825 23431 37859
rect 23673 37825 23707 37859
rect 23765 37825 23799 37859
rect 24041 37825 24075 37859
rect 24225 37825 24259 37859
rect 25053 37825 25087 37859
rect 25329 37825 25363 37859
rect 25513 37825 25547 37859
rect 25973 37825 26007 37859
rect 26433 37825 26467 37859
rect 26617 37825 26651 37859
rect 27721 37825 27755 37859
rect 28181 37825 28215 37859
rect 28825 37825 28859 37859
rect 29101 37825 29135 37859
rect 31217 37825 31251 37859
rect 10793 37757 10827 37791
rect 11713 37757 11747 37791
rect 13369 37757 13403 37791
rect 14197 37757 14231 37791
rect 14473 37757 14507 37791
rect 19901 37757 19935 37791
rect 20085 37757 20119 37791
rect 22661 37757 22695 37791
rect 25237 37757 25271 37791
rect 25697 37757 25731 37791
rect 26157 37757 26191 37791
rect 27537 37757 27571 37791
rect 27997 37757 28031 37791
rect 29377 37757 29411 37791
rect 30849 37757 30883 37791
rect 29009 37689 29043 37723
rect 13553 37621 13587 37655
rect 16497 37621 16531 37655
rect 17785 37621 17819 37655
rect 23949 37621 23983 37655
rect 28365 37621 28399 37655
rect 31033 37621 31067 37655
rect 17785 37417 17819 37451
rect 26065 37417 26099 37451
rect 27353 37417 27387 37451
rect 1685 37281 1719 37315
rect 17877 37281 17911 37315
rect 22937 37281 22971 37315
rect 26709 37281 26743 37315
rect 27997 37281 28031 37315
rect 30205 37281 30239 37315
rect 8309 37213 8343 37247
rect 8585 37213 8619 37247
rect 8677 37213 8711 37247
rect 8953 37213 8987 37247
rect 18061 37213 18095 37247
rect 18337 37213 18371 37247
rect 18521 37213 18555 37247
rect 18613 37213 18647 37247
rect 20177 37213 20211 37247
rect 20269 37213 20303 37247
rect 20453 37213 20487 37247
rect 22753 37213 22787 37247
rect 23305 37213 23339 37247
rect 23673 37213 23707 37247
rect 26433 37213 26467 37247
rect 27813 37213 27847 37247
rect 29653 37213 29687 37247
rect 29745 37213 29779 37247
rect 29929 37213 29963 37247
rect 32597 37213 32631 37247
rect 37657 37213 37691 37247
rect 1501 37145 1535 37179
rect 9229 37145 9263 37179
rect 17785 37145 17819 37179
rect 20729 37145 20763 37179
rect 22845 37145 22879 37179
rect 23489 37145 23523 37179
rect 23581 37145 23615 37179
rect 8493 37077 8527 37111
rect 10701 37077 10735 37111
rect 18245 37077 18279 37111
rect 22201 37077 22235 37111
rect 22385 37077 22419 37111
rect 23857 37077 23891 37111
rect 26525 37077 26559 37111
rect 27721 37077 27755 37111
rect 31677 37077 31711 37111
rect 32505 37077 32539 37111
rect 37841 37077 37875 37111
rect 9321 36873 9355 36907
rect 9689 36873 9723 36907
rect 20913 36873 20947 36907
rect 28089 36873 28123 36907
rect 29193 36873 29227 36907
rect 30941 36873 30975 36907
rect 31309 36873 31343 36907
rect 8769 36805 8803 36839
rect 9781 36805 9815 36839
rect 24041 36805 24075 36839
rect 7297 36737 7331 36771
rect 21097 36737 21131 36771
rect 23857 36737 23891 36771
rect 24501 36737 24535 36771
rect 24777 36737 24811 36771
rect 27721 36737 27755 36771
rect 27997 36737 28031 36771
rect 28273 36737 28307 36771
rect 29561 36737 29595 36771
rect 30849 36737 30883 36771
rect 32321 36737 32355 36771
rect 8033 36669 8067 36703
rect 9873 36669 9907 36703
rect 23673 36669 23707 36703
rect 24593 36669 24627 36703
rect 29653 36669 29687 36703
rect 29745 36669 29779 36703
rect 30665 36669 30699 36703
rect 32597 36669 32631 36703
rect 7573 36533 7607 36567
rect 24593 36533 24627 36567
rect 24961 36533 24995 36567
rect 27629 36533 27663 36567
rect 28457 36533 28491 36567
rect 34069 36533 34103 36567
rect 11805 36329 11839 36363
rect 12541 36329 12575 36363
rect 14289 36329 14323 36363
rect 15301 36329 15335 36363
rect 16497 36329 16531 36363
rect 18061 36329 18095 36363
rect 27905 36329 27939 36363
rect 32229 36329 32263 36363
rect 11989 36261 12023 36295
rect 12725 36261 12759 36295
rect 24133 36261 24167 36295
rect 32597 36261 32631 36295
rect 12633 36193 12667 36227
rect 19809 36193 19843 36227
rect 28733 36193 28767 36227
rect 33149 36193 33183 36227
rect 5733 36125 5767 36159
rect 5825 36125 5859 36159
rect 6009 36125 6043 36159
rect 9505 36125 9539 36159
rect 9781 36125 9815 36159
rect 11253 36125 11287 36159
rect 11529 36125 11563 36159
rect 11621 36125 11655 36159
rect 12111 36125 12145 36159
rect 12863 36125 12897 36159
rect 13276 36125 13310 36159
rect 13369 36125 13403 36159
rect 14289 36125 14323 36159
rect 14381 36125 14415 36159
rect 14657 36125 14691 36159
rect 14749 36125 14783 36159
rect 15301 36125 15335 36159
rect 15393 36125 15427 36159
rect 15669 36125 15703 36159
rect 15761 36125 15795 36159
rect 15945 36125 15979 36159
rect 16221 36125 16255 36159
rect 16313 36125 16347 36159
rect 16773 36125 16807 36159
rect 16866 36125 16900 36159
rect 17238 36125 17272 36159
rect 17509 36125 17543 36159
rect 17785 36125 17819 36159
rect 17877 36125 17911 36159
rect 18521 36125 18555 36159
rect 18705 36125 18739 36159
rect 20182 36125 20216 36159
rect 23581 36125 23615 36159
rect 23949 36125 23983 36159
rect 25513 36125 25547 36159
rect 25789 36125 25823 36159
rect 25881 36125 25915 36159
rect 27261 36125 27295 36159
rect 27354 36125 27388 36159
rect 27629 36125 27663 36159
rect 27767 36125 27801 36159
rect 28549 36125 28583 36159
rect 32045 36125 32079 36159
rect 33057 36125 33091 36159
rect 6285 36057 6319 36091
rect 11437 36057 11471 36091
rect 13001 36057 13035 36091
rect 13093 36057 13127 36091
rect 14565 36057 14599 36091
rect 15577 36057 15611 36091
rect 16129 36057 16163 36091
rect 17049 36057 17083 36091
rect 17141 36057 17175 36091
rect 17693 36057 17727 36091
rect 19809 36057 19843 36091
rect 19993 36057 20027 36091
rect 20085 36057 20119 36091
rect 23765 36057 23799 36091
rect 23857 36057 23891 36091
rect 25697 36057 25731 36091
rect 27537 36057 27571 36091
rect 7757 35989 7791 36023
rect 9413 35989 9447 36023
rect 9597 35989 9631 36023
rect 12173 35989 12207 36023
rect 17417 35989 17451 36023
rect 18613 35989 18647 36023
rect 26065 35989 26099 36023
rect 32965 35989 32999 36023
rect 6561 35785 6595 35819
rect 7665 35785 7699 35819
rect 13645 35785 13679 35819
rect 13921 35785 13955 35819
rect 29193 35785 29227 35819
rect 30757 35785 30791 35819
rect 9505 35717 9539 35751
rect 13277 35717 13311 35751
rect 14013 35717 14047 35751
rect 19073 35717 19107 35751
rect 21097 35717 21131 35751
rect 22201 35717 22235 35751
rect 23213 35717 23247 35751
rect 23857 35717 23891 35751
rect 25145 35717 25179 35751
rect 6745 35649 6779 35683
rect 7757 35649 7791 35683
rect 9137 35649 9171 35683
rect 9229 35649 9263 35683
rect 13093 35649 13127 35683
rect 13553 35649 13587 35683
rect 13737 35649 13771 35683
rect 14841 35649 14875 35683
rect 18889 35649 18923 35683
rect 18981 35649 19015 35683
rect 19211 35649 19245 35683
rect 21005 35649 21039 35683
rect 21189 35649 21223 35683
rect 21373 35649 21407 35683
rect 21925 35649 21959 35683
rect 22073 35649 22107 35683
rect 22290 35649 22324 35683
rect 22390 35649 22424 35683
rect 22845 35649 22879 35683
rect 22938 35649 22972 35683
rect 23121 35649 23155 35683
rect 23310 35649 23344 35683
rect 23765 35649 23799 35683
rect 23949 35649 23983 35683
rect 24133 35649 24167 35683
rect 24869 35649 24903 35683
rect 25053 35649 25087 35683
rect 25237 35649 25271 35683
rect 25697 35649 25731 35683
rect 25789 35649 25823 35683
rect 25973 35649 26007 35683
rect 26065 35649 26099 35683
rect 26157 35649 26191 35683
rect 26249 35649 26283 35683
rect 26433 35649 26467 35683
rect 26525 35649 26559 35683
rect 29653 35649 29687 35683
rect 29746 35649 29780 35683
rect 29929 35649 29963 35683
rect 30021 35649 30055 35683
rect 30118 35649 30152 35683
rect 30573 35649 30607 35683
rect 30849 35649 30883 35683
rect 31401 35649 31435 35683
rect 32965 35649 32999 35683
rect 33517 35649 33551 35683
rect 7849 35581 7883 35615
rect 8309 35581 8343 35615
rect 12909 35581 12943 35615
rect 19349 35581 19383 35615
rect 27445 35581 27479 35615
rect 27721 35581 27755 35615
rect 7297 35513 7331 35547
rect 13369 35513 13403 35547
rect 20821 35513 20855 35547
rect 22569 35513 22603 35547
rect 25421 35513 25455 35547
rect 30297 35513 30331 35547
rect 10977 35445 11011 35479
rect 18705 35445 18739 35479
rect 23489 35445 23523 35479
rect 23581 35445 23615 35479
rect 25513 35445 25547 35479
rect 26709 35445 26743 35479
rect 30389 35445 30423 35479
rect 31217 35445 31251 35479
rect 32873 35445 32907 35479
rect 33333 35445 33367 35479
rect 9505 35241 9539 35275
rect 17509 35241 17543 35275
rect 28181 35241 28215 35275
rect 28089 35173 28123 35207
rect 9965 35105 9999 35139
rect 10057 35105 10091 35139
rect 23581 35105 23615 35139
rect 23673 35105 23707 35139
rect 26065 35105 26099 35139
rect 27537 35105 27571 35139
rect 30941 35105 30975 35139
rect 32689 35105 32723 35139
rect 32965 35105 32999 35139
rect 6653 35037 6687 35071
rect 6745 35037 6779 35071
rect 6929 35037 6963 35071
rect 9873 35037 9907 35071
rect 17325 35037 17359 35071
rect 23305 35037 23339 35071
rect 23489 35037 23523 35071
rect 23765 35037 23799 35071
rect 25329 35037 25363 35071
rect 25513 35037 25547 35071
rect 25605 35037 25639 35071
rect 25697 35037 25731 35071
rect 26341 35037 26375 35071
rect 26433 35037 26467 35071
rect 26525 35037 26559 35071
rect 26709 35037 26743 35071
rect 27721 35037 27755 35071
rect 28365 35037 28399 35071
rect 28917 35037 28951 35071
rect 30389 35037 30423 35071
rect 30481 35037 30515 35071
rect 30665 35037 30699 35071
rect 7205 34969 7239 35003
rect 8677 34901 8711 34935
rect 23949 34901 23983 34935
rect 25973 34901 26007 34935
rect 27629 34901 27663 34935
rect 28825 34901 28859 34935
rect 32413 34901 32447 34935
rect 34437 34901 34471 34935
rect 7665 34697 7699 34731
rect 7941 34697 7975 34731
rect 16865 34697 16899 34731
rect 31217 34697 31251 34731
rect 33333 34697 33367 34731
rect 33701 34697 33735 34731
rect 11805 34629 11839 34663
rect 17233 34629 17267 34663
rect 21005 34629 21039 34663
rect 21221 34629 21255 34663
rect 22201 34629 22235 34663
rect 23581 34629 23615 34663
rect 5641 34561 5675 34595
rect 7849 34561 7883 34595
rect 8309 34561 8343 34595
rect 11708 34561 11742 34595
rect 11897 34561 11931 34595
rect 12080 34561 12114 34595
rect 12173 34561 12207 34595
rect 17141 34561 17175 34595
rect 21925 34561 21959 34595
rect 22018 34561 22052 34595
rect 22293 34561 22327 34595
rect 22390 34561 22424 34595
rect 23397 34561 23431 34595
rect 23673 34561 23707 34595
rect 23765 34561 23799 34595
rect 28641 34561 28675 34595
rect 31585 34561 31619 34595
rect 37565 34561 37599 34595
rect 8401 34493 8435 34527
rect 8585 34493 8619 34527
rect 31677 34493 31711 34527
rect 31769 34493 31803 34527
rect 33057 34493 33091 34527
rect 33241 34493 33275 34527
rect 37841 34493 37875 34527
rect 21373 34425 21407 34459
rect 5457 34357 5491 34391
rect 11529 34357 11563 34391
rect 16865 34357 16899 34391
rect 16957 34357 16991 34391
rect 17049 34357 17083 34391
rect 21189 34357 21223 34391
rect 22569 34357 22603 34391
rect 23949 34357 23983 34391
rect 28898 34357 28932 34391
rect 30389 34357 30423 34391
rect 14841 34153 14875 34187
rect 15117 34153 15151 34187
rect 16681 34153 16715 34187
rect 28089 34153 28123 34187
rect 11621 34085 11655 34119
rect 15945 34085 15979 34119
rect 19441 34085 19475 34119
rect 19901 34085 19935 34119
rect 26065 34085 26099 34119
rect 28457 34085 28491 34119
rect 31125 34085 31159 34119
rect 34069 34085 34103 34119
rect 13185 34017 13219 34051
rect 13737 34017 13771 34051
rect 14749 34017 14783 34051
rect 15393 34017 15427 34051
rect 16865 34017 16899 34051
rect 29101 34017 29135 34051
rect 34989 34017 35023 34051
rect 4721 33949 4755 33983
rect 4813 33949 4847 33983
rect 4997 33949 5031 33983
rect 7297 33949 7331 33983
rect 8585 33949 8619 33983
rect 9505 33949 9539 33983
rect 9873 33949 9907 33983
rect 11621 33949 11655 33983
rect 11805 33949 11839 33983
rect 11897 33949 11931 33983
rect 13461 33949 13495 33983
rect 14381 33949 14415 33983
rect 14565 33949 14599 33983
rect 14657 33949 14691 33983
rect 16037 33949 16071 33983
rect 16221 33949 16255 33983
rect 16313 33949 16347 33983
rect 16405 33949 16439 33983
rect 17049 33949 17083 33983
rect 17233 33949 17267 33983
rect 17417 33949 17451 33983
rect 17693 33949 17727 33983
rect 17786 33949 17820 33983
rect 18158 33949 18192 33983
rect 18429 33949 18463 33983
rect 18705 33949 18739 33983
rect 18797 33949 18831 33983
rect 19257 33949 19291 33983
rect 19533 33949 19567 33983
rect 20085 33949 20119 33983
rect 20269 33949 20303 33983
rect 20453 33949 20487 33983
rect 20821 33949 20855 33983
rect 21925 33949 21959 33983
rect 22109 33949 22143 33983
rect 22569 33949 22603 33983
rect 22661 33949 22695 33983
rect 22845 33949 22879 33983
rect 22937 33949 22971 33983
rect 23213 33949 23247 33983
rect 23306 33949 23340 33983
rect 23489 33949 23523 33983
rect 23581 33949 23615 33983
rect 23719 33949 23753 33983
rect 25605 33949 25639 33983
rect 25697 33949 25731 33983
rect 25881 33949 25915 33983
rect 25973 33949 26007 33983
rect 26249 33949 26283 33983
rect 26341 33949 26375 33983
rect 26617 33949 26651 33983
rect 27261 33949 27295 33983
rect 27905 33949 27939 33983
rect 30481 33949 30515 33983
rect 30574 33949 30608 33983
rect 30849 33949 30883 33983
rect 30946 33949 30980 33983
rect 31493 33949 31527 33983
rect 31769 33949 31803 33983
rect 33885 33949 33919 33983
rect 34345 33949 34379 33983
rect 34437 33949 34471 33983
rect 34713 33949 34747 33983
rect 5273 33881 5307 33915
rect 15577 33881 15611 33915
rect 17969 33881 18003 33915
rect 18061 33881 18095 33915
rect 18613 33881 18647 33915
rect 20177 33881 20211 33915
rect 26433 33881 26467 33915
rect 28917 33881 28951 33915
rect 30757 33881 30791 33915
rect 36737 33881 36771 33915
rect 6745 33813 6779 33847
rect 7205 33813 7239 33847
rect 8677 33813 8711 33847
rect 8953 33813 8987 33847
rect 9689 33813 9723 33847
rect 13369 33813 13403 33847
rect 13553 33813 13587 33847
rect 15669 33813 15703 33847
rect 15761 33813 15795 33847
rect 17141 33813 17175 33847
rect 18337 33813 18371 33847
rect 18981 33813 19015 33847
rect 19533 33813 19567 33847
rect 23121 33813 23155 33847
rect 23857 33813 23891 33847
rect 25421 33813 25455 33847
rect 27169 33813 27203 33847
rect 28825 33813 28859 33847
rect 31585 33813 31619 33847
rect 31953 33813 31987 33847
rect 5457 33609 5491 33643
rect 5825 33609 5859 33643
rect 14381 33609 14415 33643
rect 14565 33609 14599 33643
rect 17601 33609 17635 33643
rect 21097 33609 21131 33643
rect 21281 33609 21315 33643
rect 33333 33609 33367 33643
rect 33793 33609 33827 33643
rect 34161 33609 34195 33643
rect 34621 33609 34655 33643
rect 36921 33609 36955 33643
rect 9229 33541 9263 33575
rect 14289 33541 14323 33575
rect 17233 33541 17267 33575
rect 20821 33541 20855 33575
rect 21465 33541 21499 33575
rect 25237 33541 25271 33575
rect 17463 33507 17497 33541
rect 7021 33473 7055 33507
rect 8953 33473 8987 33507
rect 14197 33473 14231 33507
rect 19708 33473 19742 33507
rect 19901 33473 19935 33507
rect 20269 33473 20303 33507
rect 20361 33473 20395 33507
rect 20637 33473 20671 33507
rect 20729 33473 20763 33507
rect 20913 33473 20947 33507
rect 21833 33473 21867 33507
rect 22017 33473 22051 33507
rect 23765 33473 23799 33507
rect 23857 33473 23891 33507
rect 26617 33473 26651 33507
rect 26985 33473 27019 33507
rect 33425 33473 33459 33507
rect 34253 33473 34287 33507
rect 34713 33473 34747 33507
rect 36737 33473 36771 33507
rect 5917 33405 5951 33439
rect 6101 33405 6135 33439
rect 7297 33405 7331 33439
rect 8769 33405 8803 33439
rect 14013 33405 14047 33439
rect 19073 33405 19107 33439
rect 23489 33405 23523 33439
rect 23581 33405 23615 33439
rect 27261 33405 27295 33439
rect 29009 33405 29043 33439
rect 33241 33405 33275 33439
rect 34069 33405 34103 33439
rect 21833 33337 21867 33371
rect 24869 33337 24903 33371
rect 26801 33337 26835 33371
rect 10701 33269 10735 33303
rect 17417 33269 17451 33303
rect 21281 33269 21315 33303
rect 24041 33269 24075 33303
rect 25237 33269 25271 33303
rect 25421 33269 25455 33303
rect 34897 33269 34931 33303
rect 7665 33065 7699 33099
rect 10149 33065 10183 33099
rect 18613 33065 18647 33099
rect 26617 33065 26651 33099
rect 19809 32997 19843 33031
rect 6101 32929 6135 32963
rect 6745 32929 6779 32963
rect 6837 32929 6871 32963
rect 8125 32929 8159 32963
rect 8401 32929 8435 32963
rect 9597 32929 9631 32963
rect 19629 32929 19663 32963
rect 22293 32929 22327 32963
rect 27169 32929 27203 32963
rect 34989 32929 35023 32963
rect 4077 32861 4111 32895
rect 4169 32861 4203 32895
rect 4353 32861 4387 32895
rect 6653 32861 6687 32895
rect 7849 32861 7883 32895
rect 7941 32861 7975 32895
rect 8217 32861 8251 32895
rect 8493 32861 8527 32895
rect 9781 32861 9815 32895
rect 11713 32861 11747 32895
rect 11851 32861 11885 32895
rect 12178 32861 12212 32895
rect 16221 32861 16255 32895
rect 16865 32861 16899 32895
rect 18337 32861 18371 32895
rect 18705 32861 18739 32895
rect 19901 32861 19935 32895
rect 20177 32861 20211 32895
rect 20453 32861 20487 32895
rect 20545 32861 20579 32895
rect 21465 32861 21499 32895
rect 22109 32861 22143 32895
rect 23397 32861 23431 32895
rect 27537 32861 27571 32895
rect 30389 32861 30423 32895
rect 30941 32861 30975 32895
rect 31217 32861 31251 32895
rect 34345 32861 34379 32895
rect 34437 32861 34471 32895
rect 34713 32861 34747 32895
rect 4629 32793 4663 32827
rect 11989 32793 12023 32827
rect 12081 32793 12115 32827
rect 18429 32793 18463 32827
rect 18797 32793 18831 32827
rect 19625 32793 19659 32827
rect 20361 32793 20395 32827
rect 23213 32793 23247 32827
rect 27813 32793 27847 32827
rect 31493 32793 31527 32827
rect 36737 32793 36771 32827
rect 6285 32725 6319 32759
rect 9689 32725 9723 32759
rect 12357 32725 12391 32759
rect 16405 32725 16439 32759
rect 20729 32725 20763 32759
rect 23581 32725 23615 32759
rect 26985 32725 27019 32759
rect 27077 32725 27111 32759
rect 29285 32725 29319 32759
rect 30205 32725 30239 32759
rect 31125 32725 31159 32759
rect 32965 32725 32999 32759
rect 4997 32521 5031 32555
rect 12081 32521 12115 32555
rect 16865 32521 16899 32555
rect 17693 32521 17727 32555
rect 27813 32521 27847 32555
rect 29009 32521 29043 32555
rect 31401 32521 31435 32555
rect 36001 32521 36035 32555
rect 11805 32453 11839 32487
rect 12265 32453 12299 32487
rect 12449 32453 12483 32487
rect 16681 32453 16715 32487
rect 17325 32453 17359 32487
rect 17509 32453 17543 32487
rect 23121 32453 23155 32487
rect 23213 32453 23247 32487
rect 23949 32453 23983 32487
rect 5181 32385 5215 32419
rect 11529 32385 11563 32419
rect 11713 32385 11747 32419
rect 11897 32385 11931 32419
rect 18429 32385 18463 32419
rect 18613 32385 18647 32419
rect 18705 32385 18739 32419
rect 18889 32385 18923 32419
rect 18981 32385 19015 32419
rect 21281 32385 21315 32419
rect 21925 32385 21959 32419
rect 23029 32385 23063 32419
rect 23397 32385 23431 32419
rect 23765 32385 23799 32419
rect 24041 32385 24075 32419
rect 24133 32385 24167 32419
rect 27905 32385 27939 32419
rect 28549 32385 28583 32419
rect 29193 32385 29227 32419
rect 30757 32385 30791 32419
rect 30849 32385 30883 32419
rect 31493 32385 31527 32419
rect 32413 32385 32447 32419
rect 33149 32385 33183 32419
rect 33425 32385 33459 32419
rect 35633 32385 35667 32419
rect 35817 32385 35851 32419
rect 28273 32317 28307 32351
rect 28457 32317 28491 32351
rect 30665 32317 30699 32351
rect 32689 32317 32723 32351
rect 12633 32249 12667 32283
rect 17049 32249 17083 32283
rect 28917 32249 28951 32283
rect 31217 32249 31251 32283
rect 32873 32249 32907 32283
rect 16865 32181 16899 32215
rect 17509 32181 17543 32215
rect 19993 32181 20027 32215
rect 22201 32181 22235 32215
rect 22845 32181 22879 32215
rect 24317 32181 24351 32215
rect 4524 31977 4558 32011
rect 7297 31977 7331 32011
rect 19073 31977 19107 32011
rect 24041 31977 24075 32011
rect 24961 31909 24995 31943
rect 25237 31909 25271 31943
rect 26801 31909 26835 31943
rect 30205 31909 30239 31943
rect 6285 31841 6319 31875
rect 6653 31841 6687 31875
rect 7205 31841 7239 31875
rect 3985 31773 4019 31807
rect 4077 31773 4111 31807
rect 4261 31773 4295 31807
rect 7481 31773 7515 31807
rect 7573 31773 7607 31807
rect 7665 31773 7699 31807
rect 7849 31773 7883 31807
rect 8125 31773 8159 31807
rect 8493 31773 8527 31807
rect 9229 31773 9263 31807
rect 9321 31773 9355 31807
rect 9505 31773 9539 31807
rect 13645 31773 13679 31807
rect 18889 31773 18923 31807
rect 19073 31773 19107 31807
rect 21281 31773 21315 31807
rect 21925 31773 21959 31807
rect 22018 31773 22052 31807
rect 22201 31773 22235 31807
rect 22293 31773 22327 31807
rect 22390 31773 22424 31807
rect 22661 31773 22695 31807
rect 22809 31773 22843 31807
rect 23126 31773 23160 31807
rect 23397 31773 23431 31807
rect 23490 31773 23524 31807
rect 23673 31773 23707 31807
rect 23903 31773 23937 31807
rect 24409 31773 24443 31807
rect 24777 31773 24811 31807
rect 25145 31773 25179 31807
rect 25329 31773 25363 31807
rect 25421 31773 25455 31807
rect 26157 31773 26191 31807
rect 26249 31773 26283 31807
rect 26525 31773 26559 31807
rect 26985 31773 27019 31807
rect 27997 31773 28031 31807
rect 28273 31773 28307 31807
rect 29561 31773 29595 31807
rect 29654 31773 29688 31807
rect 29837 31773 29871 31807
rect 29929 31773 29963 31807
rect 30026 31773 30060 31807
rect 30481 31773 30515 31807
rect 31493 31773 31527 31807
rect 31769 31773 31803 31807
rect 34897 31773 34931 31807
rect 34989 31773 35023 31807
rect 35449 31773 35483 31807
rect 9781 31705 9815 31739
rect 13093 31705 13127 31739
rect 13277 31705 13311 31739
rect 22937 31705 22971 31739
rect 23029 31705 23063 31739
rect 23765 31705 23799 31739
rect 24593 31705 24627 31739
rect 24685 31705 24719 31739
rect 26341 31705 26375 31739
rect 31585 31705 31619 31739
rect 35081 31705 35115 31739
rect 8033 31637 8067 31671
rect 8309 31637 8343 31671
rect 11253 31637 11287 31671
rect 13369 31637 13403 31671
rect 13461 31637 13495 31671
rect 18705 31637 18739 31671
rect 19993 31637 20027 31671
rect 22569 31637 22603 31671
rect 23305 31637 23339 31671
rect 25605 31637 25639 31671
rect 25973 31637 26007 31671
rect 27905 31637 27939 31671
rect 28089 31637 28123 31671
rect 30389 31637 30423 31671
rect 31953 31637 31987 31671
rect 34805 31637 34839 31671
rect 35265 31637 35299 31671
rect 9873 31433 9907 31467
rect 10149 31433 10183 31467
rect 13461 31433 13495 31467
rect 17325 31433 17359 31467
rect 18705 31433 18739 31467
rect 22109 31433 22143 31467
rect 22201 31433 22235 31467
rect 22385 31433 22419 31467
rect 8125 31365 8159 31399
rect 11713 31365 11747 31399
rect 14749 31365 14783 31399
rect 16129 31365 16163 31399
rect 23397 31365 23431 31399
rect 25145 31365 25179 31399
rect 27997 31365 28031 31399
rect 10057 31297 10091 31331
rect 10517 31297 10551 31331
rect 11529 31297 11563 31331
rect 11805 31297 11839 31331
rect 11897 31297 11931 31331
rect 15485 31297 15519 31331
rect 15669 31297 15703 31331
rect 15945 31297 15979 31331
rect 16221 31297 16255 31331
rect 16313 31297 16347 31331
rect 16670 31297 16704 31331
rect 16829 31297 16863 31331
rect 16957 31297 16991 31331
rect 17049 31297 17083 31331
rect 17165 31297 17199 31331
rect 17417 31297 17451 31331
rect 17601 31297 17635 31331
rect 17693 31297 17727 31331
rect 17785 31297 17819 31331
rect 18521 31297 18555 31331
rect 18797 31297 18831 31331
rect 19257 31297 19291 31331
rect 19533 31297 19567 31331
rect 19717 31297 19751 31331
rect 20545 31297 20579 31331
rect 20637 31297 20671 31331
rect 20821 31297 20855 31331
rect 20913 31297 20947 31331
rect 21373 31297 21407 31331
rect 21465 31297 21499 31331
rect 21833 31297 21867 31331
rect 22017 31297 22051 31331
rect 22845 31297 22879 31331
rect 23029 31297 23063 31331
rect 23305 31297 23339 31331
rect 25421 31297 25455 31331
rect 25605 31297 25639 31331
rect 26341 31297 26375 31331
rect 26985 31297 27019 31331
rect 27169 31297 27203 31331
rect 27261 31297 27295 31331
rect 27353 31297 27387 31331
rect 29653 31297 29687 31331
rect 29929 31297 29963 31331
rect 32413 31297 32447 31331
rect 34437 31297 34471 31331
rect 34529 31297 34563 31331
rect 7849 31229 7883 31263
rect 10609 31229 10643 31263
rect 10793 31229 10827 31263
rect 15393 31229 15427 31263
rect 15853 31229 15887 31263
rect 21005 31229 21039 31263
rect 21189 31229 21223 31263
rect 21281 31229 21315 31263
rect 22937 31229 22971 31263
rect 23121 31229 23155 31263
rect 26065 31229 26099 31263
rect 27721 31229 27755 31263
rect 30205 31229 30239 31263
rect 31953 31229 31987 31263
rect 34161 31229 34195 31263
rect 34805 31229 34839 31263
rect 36553 31229 36587 31263
rect 9597 31161 9631 31195
rect 26709 31161 26743 31195
rect 29837 31161 29871 31195
rect 12081 31093 12115 31127
rect 16497 31093 16531 31127
rect 17969 31093 18003 31127
rect 18337 31093 18371 31127
rect 20361 31093 20395 31127
rect 22661 31093 22695 31127
rect 27629 31093 27663 31127
rect 29469 31093 29503 31127
rect 8953 30889 8987 30923
rect 14473 30889 14507 30923
rect 16497 30889 16531 30923
rect 21281 30889 21315 30923
rect 24501 30889 24535 30923
rect 24869 30889 24903 30923
rect 26617 30889 26651 30923
rect 28089 30889 28123 30923
rect 30113 30889 30147 30923
rect 34069 30889 34103 30923
rect 35449 30889 35483 30923
rect 13369 30821 13403 30855
rect 20361 30821 20395 30855
rect 20729 30821 20763 30855
rect 21741 30821 21775 30855
rect 33793 30821 33827 30855
rect 7665 30753 7699 30787
rect 8401 30753 8435 30787
rect 9413 30753 9447 30787
rect 9505 30753 9539 30787
rect 13921 30753 13955 30787
rect 14565 30753 14599 30787
rect 24593 30753 24627 30787
rect 28641 30753 28675 30787
rect 30665 30753 30699 30787
rect 33149 30753 33183 30787
rect 34805 30753 34839 30787
rect 4537 30685 4571 30719
rect 5641 30685 5675 30719
rect 5733 30685 5767 30719
rect 5917 30685 5951 30719
rect 8217 30685 8251 30719
rect 14381 30685 14415 30719
rect 14657 30685 14691 30719
rect 14841 30685 14875 30719
rect 16313 30685 16347 30719
rect 16589 30685 16623 30719
rect 16682 30685 16716 30719
rect 16865 30685 16899 30719
rect 17095 30685 17129 30719
rect 19073 30685 19107 30719
rect 19533 30685 19567 30719
rect 20269 30685 20303 30719
rect 21097 30685 21131 30719
rect 21373 30685 21407 30719
rect 24501 30685 24535 30719
rect 26065 30685 26099 30719
rect 26157 30685 26191 30719
rect 26341 30685 26375 30719
rect 26433 30685 26467 30719
rect 30481 30685 30515 30719
rect 33425 30685 33459 30719
rect 33885 30685 33919 30719
rect 6193 30617 6227 30651
rect 13737 30617 13771 30651
rect 16129 30617 16163 30651
rect 16957 30617 16991 30651
rect 21005 30617 21039 30651
rect 21557 30617 21591 30651
rect 28549 30617 28583 30651
rect 30941 30617 30975 30651
rect 34989 30617 35023 30651
rect 4445 30549 4479 30583
rect 7849 30549 7883 30583
rect 8309 30549 8343 30583
rect 9321 30549 9355 30583
rect 13553 30549 13587 30583
rect 13645 30549 13679 30583
rect 14105 30549 14139 30583
rect 17233 30549 17267 30583
rect 17785 30549 17819 30583
rect 20913 30549 20947 30583
rect 28457 30549 28491 30583
rect 30573 30549 30607 30583
rect 32229 30549 32263 30583
rect 33333 30549 33367 30583
rect 35081 30549 35115 30583
rect 6009 30345 6043 30379
rect 6469 30345 6503 30379
rect 20269 30345 20303 30379
rect 29101 30345 29135 30379
rect 7389 30277 7423 30311
rect 13001 30277 13035 30311
rect 14749 30277 14783 30311
rect 19901 30277 19935 30311
rect 20085 30277 20119 30311
rect 20453 30277 20487 30311
rect 20637 30277 20671 30311
rect 23397 30277 23431 30311
rect 6653 30209 6687 30243
rect 7665 30209 7699 30243
rect 7757 30209 7791 30243
rect 7849 30209 7883 30243
rect 8033 30209 8067 30243
rect 8585 30209 8619 30243
rect 11621 30209 11655 30243
rect 11714 30209 11748 30243
rect 11897 30209 11931 30243
rect 11989 30209 12023 30243
rect 12127 30209 12161 30243
rect 17693 30209 17727 30243
rect 18429 30209 18463 30243
rect 18521 30209 18555 30243
rect 18613 30209 18647 30243
rect 18797 30209 18831 30243
rect 25697 30209 25731 30243
rect 25881 30209 25915 30243
rect 25973 30209 26007 30243
rect 26065 30209 26099 30243
rect 30389 30209 30423 30243
rect 32137 30209 32171 30243
rect 32321 30209 32355 30243
rect 32413 30209 32447 30243
rect 32505 30209 32539 30243
rect 4261 30141 4295 30175
rect 4537 30141 4571 30175
rect 6745 30141 6779 30175
rect 17785 30141 17819 30175
rect 25145 30141 25179 30175
rect 7481 30073 7515 30107
rect 18061 30073 18095 30107
rect 8677 30005 8711 30039
rect 12265 30005 12299 30039
rect 17877 30005 17911 30039
rect 18153 30005 18187 30039
rect 20085 30005 20119 30039
rect 20637 30005 20671 30039
rect 20821 30005 20855 30039
rect 26249 30005 26283 30039
rect 32781 30005 32815 30039
rect 10701 29801 10735 29835
rect 12541 29801 12575 29835
rect 15761 29801 15795 29835
rect 16681 29801 16715 29835
rect 24593 29801 24627 29835
rect 8493 29733 8527 29767
rect 13737 29733 13771 29767
rect 14105 29733 14139 29767
rect 14381 29733 14415 29767
rect 15117 29733 15151 29767
rect 18889 29733 18923 29767
rect 20637 29733 20671 29767
rect 6101 29665 6135 29699
rect 9229 29665 9263 29699
rect 14473 29665 14507 29699
rect 24685 29665 24719 29699
rect 26249 29665 26283 29699
rect 27629 29665 27663 29699
rect 33977 29665 34011 29699
rect 36829 29665 36863 29699
rect 4169 29597 4203 29631
rect 5917 29597 5951 29631
rect 8309 29597 8343 29631
rect 8585 29597 8619 29631
rect 8677 29597 8711 29631
rect 8953 29597 8987 29631
rect 12725 29597 12759 29631
rect 12909 29597 12943 29631
rect 13461 29597 13495 29631
rect 13553 29597 13587 29631
rect 13829 29597 13863 29631
rect 14289 29597 14323 29631
rect 14565 29597 14599 29631
rect 14749 29597 14783 29631
rect 15301 29597 15335 29631
rect 15393 29597 15427 29631
rect 15485 29597 15519 29631
rect 15669 29597 15703 29631
rect 15945 29597 15979 29631
rect 16129 29597 16163 29631
rect 16313 29597 16347 29631
rect 18245 29597 18279 29631
rect 18337 29597 18371 29631
rect 18521 29597 18555 29631
rect 18613 29597 18647 29631
rect 18705 29597 18739 29631
rect 20913 29597 20947 29631
rect 21005 29597 21039 29631
rect 22932 29597 22966 29631
rect 23121 29597 23155 29631
rect 23249 29597 23283 29631
rect 23397 29597 23431 29631
rect 23765 29597 23799 29631
rect 24041 29597 24075 29631
rect 24777 29597 24811 29631
rect 25789 29597 25823 29631
rect 25881 29597 25915 29631
rect 25973 29597 26007 29631
rect 26157 29597 26191 29631
rect 26433 29597 26467 29631
rect 26525 29597 26559 29631
rect 26709 29597 26743 29631
rect 26801 29597 26835 29631
rect 27353 29597 27387 29631
rect 27445 29597 27479 29631
rect 28549 29597 28583 29631
rect 29377 29597 29411 29631
rect 29837 29597 29871 29631
rect 29929 29597 29963 29631
rect 30021 29597 30055 29631
rect 30205 29597 30239 29631
rect 30297 29597 30331 29631
rect 30390 29597 30424 29631
rect 30573 29597 30607 29631
rect 30803 29597 30837 29631
rect 31217 29597 31251 29631
rect 34161 29597 34195 29631
rect 34805 29597 34839 29631
rect 5825 29529 5859 29563
rect 16037 29529 16071 29563
rect 17233 29529 17267 29563
rect 23029 29529 23063 29563
rect 30665 29529 30699 29563
rect 32965 29529 32999 29563
rect 35081 29529 35115 29563
rect 4077 29461 4111 29495
rect 5457 29461 5491 29495
rect 13277 29461 13311 29495
rect 16865 29461 16899 29495
rect 16957 29461 16991 29495
rect 17049 29461 17083 29495
rect 20821 29461 20855 29495
rect 21189 29461 21223 29495
rect 22753 29461 22787 29495
rect 23581 29461 23615 29495
rect 23949 29461 23983 29495
rect 24409 29461 24443 29495
rect 25513 29461 25547 29495
rect 27813 29461 27847 29495
rect 27905 29461 27939 29495
rect 28273 29461 28307 29495
rect 28365 29461 28399 29495
rect 29285 29461 29319 29495
rect 29561 29461 29595 29495
rect 30941 29461 30975 29495
rect 34069 29461 34103 29495
rect 34529 29461 34563 29495
rect 8769 29257 8803 29291
rect 9137 29257 9171 29291
rect 18889 29257 18923 29291
rect 29009 29257 29043 29291
rect 31585 29257 31619 29291
rect 34989 29257 35023 29291
rect 7021 29189 7055 29223
rect 11345 29189 11379 29223
rect 20913 29189 20947 29223
rect 23673 29189 23707 29223
rect 26065 29189 26099 29223
rect 27537 29189 27571 29223
rect 3893 29121 3927 29155
rect 6929 29121 6963 29155
rect 7113 29121 7147 29155
rect 7297 29121 7331 29155
rect 7665 29121 7699 29155
rect 13093 29121 13127 29155
rect 13277 29121 13311 29155
rect 18521 29121 18555 29155
rect 18705 29121 18739 29155
rect 20729 29121 20763 29155
rect 21005 29121 21039 29155
rect 21097 29121 21131 29155
rect 21833 29121 21867 29155
rect 21981 29121 22015 29155
rect 22109 29121 22143 29155
rect 22201 29121 22235 29155
rect 22298 29121 22332 29155
rect 22569 29121 22603 29155
rect 22845 29121 22879 29155
rect 23029 29121 23063 29155
rect 23489 29121 23523 29155
rect 23765 29121 23799 29155
rect 23857 29121 23891 29155
rect 25513 29121 25547 29155
rect 25605 29121 25639 29155
rect 25789 29121 25823 29155
rect 25881 29121 25915 29155
rect 26157 29121 26191 29155
rect 26341 29121 26375 29155
rect 26433 29121 26467 29155
rect 26525 29121 26559 29155
rect 27261 29121 27295 29155
rect 29193 29121 29227 29155
rect 31493 29121 31527 29155
rect 31769 29121 31803 29155
rect 31953 29121 31987 29155
rect 32137 29121 32171 29155
rect 32321 29121 32355 29155
rect 32413 29121 32447 29155
rect 32506 29143 32540 29177
rect 33057 29121 33091 29155
rect 34621 29121 34655 29155
rect 35081 29121 35115 29155
rect 36645 29121 36679 29155
rect 36829 29121 36863 29155
rect 5917 29053 5951 29087
rect 8309 29053 8343 29087
rect 9229 29053 9263 29087
rect 9413 29053 9447 29087
rect 22753 29053 22787 29087
rect 30941 29053 30975 29087
rect 9873 28985 9907 29019
rect 12909 28985 12943 29019
rect 22477 28985 22511 29019
rect 22937 28985 22971 29019
rect 26801 28985 26835 29019
rect 32781 28985 32815 29019
rect 34805 28985 34839 29019
rect 37013 28985 37047 29019
rect 4156 28917 4190 28951
rect 6745 28917 6779 28951
rect 18613 28917 18647 28951
rect 21281 28917 21315 28951
rect 23213 28917 23247 28951
rect 24041 28917 24075 28951
rect 29450 28917 29484 28951
rect 32873 28917 32907 28951
rect 4537 28713 4571 28747
rect 7941 28713 7975 28747
rect 25789 28713 25823 28747
rect 29285 28713 29319 28747
rect 6009 28577 6043 28611
rect 6193 28577 6227 28611
rect 6469 28577 6503 28611
rect 30021 28577 30055 28611
rect 30113 28577 30147 28611
rect 32045 28577 32079 28611
rect 33885 28577 33919 28611
rect 34069 28577 34103 28611
rect 36461 28577 36495 28611
rect 4353 28509 4387 28543
rect 4721 28509 4755 28543
rect 6101 28509 6135 28543
rect 8309 28509 8343 28543
rect 9965 28509 9999 28543
rect 10057 28509 10091 28543
rect 10241 28509 10275 28543
rect 16129 28509 16163 28543
rect 16313 28509 16347 28543
rect 16497 28509 16531 28543
rect 19717 28509 19751 28543
rect 19809 28509 19843 28543
rect 20085 28509 20119 28543
rect 20821 28509 20855 28543
rect 22477 28509 22511 28543
rect 24593 28509 24627 28543
rect 24685 28509 24719 28543
rect 24961 28509 24995 28543
rect 25973 28509 26007 28543
rect 26065 28509 26099 28543
rect 26341 28509 26375 28543
rect 29101 28509 29135 28543
rect 30389 28509 30423 28543
rect 30482 28509 30516 28543
rect 30757 28509 30791 28543
rect 30854 28509 30888 28543
rect 31309 28509 31343 28543
rect 31585 28509 31619 28543
rect 31769 28509 31803 28543
rect 34713 28509 34747 28543
rect 10517 28441 10551 28475
rect 16405 28441 16439 28475
rect 19901 28441 19935 28475
rect 24777 28441 24811 28475
rect 26157 28441 26191 28475
rect 30665 28441 30699 28475
rect 34989 28441 35023 28475
rect 4261 28373 4295 28407
rect 8217 28373 8251 28407
rect 11989 28373 12023 28407
rect 16681 28373 16715 28407
rect 19533 28373 19567 28407
rect 24409 28373 24443 28407
rect 29561 28373 29595 28407
rect 29929 28373 29963 28407
rect 31033 28373 31067 28407
rect 31125 28373 31159 28407
rect 31493 28373 31527 28407
rect 33517 28373 33551 28407
rect 34161 28373 34195 28407
rect 34529 28373 34563 28407
rect 6837 28169 6871 28203
rect 10609 28169 10643 28203
rect 11529 28169 11563 28203
rect 11897 28169 11931 28203
rect 13737 28169 13771 28203
rect 13921 28169 13955 28203
rect 14841 28169 14875 28203
rect 23121 28169 23155 28203
rect 23857 28169 23891 28203
rect 31861 28169 31895 28203
rect 32597 28169 32631 28203
rect 32965 28169 32999 28203
rect 34437 28169 34471 28203
rect 34897 28169 34931 28203
rect 4353 28101 4387 28135
rect 12633 28101 12667 28135
rect 17049 28101 17083 28135
rect 19073 28101 19107 28135
rect 19273 28101 19307 28135
rect 4077 28033 4111 28067
rect 6745 28033 6779 28067
rect 7665 28033 7699 28067
rect 9965 28033 9999 28067
rect 10793 28033 10827 28067
rect 12469 28033 12503 28067
rect 12725 28033 12759 28067
rect 12817 28033 12851 28067
rect 13829 28033 13863 28067
rect 14933 28033 14967 28067
rect 16681 28033 16715 28067
rect 16774 28033 16808 28067
rect 16957 28033 16991 28067
rect 17187 28033 17221 28067
rect 19625 28033 19659 28067
rect 19911 28033 19945 28067
rect 20085 28033 20119 28067
rect 20637 28033 20671 28067
rect 20821 28033 20855 28067
rect 20914 28033 20948 28067
rect 21097 28033 21131 28067
rect 21189 28033 21223 28067
rect 21286 28033 21320 28067
rect 22477 28033 22511 28067
rect 22845 28033 22879 28067
rect 23305 28033 23339 28067
rect 23397 28033 23431 28067
rect 23489 28033 23523 28067
rect 23673 28033 23707 28067
rect 23765 28033 23799 28067
rect 24133 28033 24167 28067
rect 31953 28033 31987 28067
rect 32505 28033 32539 28067
rect 34253 28033 34287 28067
rect 34989 28033 35023 28067
rect 37381 28033 37415 28067
rect 5825 27965 5859 27999
rect 7021 27965 7055 27999
rect 7941 27965 7975 27999
rect 9413 27965 9447 27999
rect 10057 27965 10091 27999
rect 10149 27965 10183 27999
rect 11989 27965 12023 27999
rect 12081 27965 12115 27999
rect 13553 27965 13587 27999
rect 19809 27965 19843 27999
rect 20177 27965 20211 27999
rect 20361 27965 20395 27999
rect 20453 27965 20487 27999
rect 20545 27965 20579 27999
rect 21925 27965 21959 27999
rect 22293 27965 22327 27999
rect 22753 27965 22787 27999
rect 32413 27965 32447 27999
rect 14105 27897 14139 27931
rect 14565 27897 14599 27931
rect 14657 27897 14691 27931
rect 19441 27897 19475 27931
rect 19717 27897 19751 27931
rect 21465 27897 21499 27931
rect 24041 27897 24075 27931
rect 6377 27829 6411 27863
rect 9597 27829 9631 27863
rect 13001 27829 13035 27863
rect 14197 27829 14231 27863
rect 14473 27829 14507 27863
rect 17325 27829 17359 27863
rect 19257 27829 19291 27863
rect 24225 27829 24259 27863
rect 24501 27829 24535 27863
rect 37565 27829 37599 27863
rect 4629 27625 4663 27659
rect 8309 27625 8343 27659
rect 14657 27625 14691 27659
rect 16037 27625 16071 27659
rect 23765 27625 23799 27659
rect 14105 27557 14139 27591
rect 33793 27557 33827 27591
rect 12081 27489 12115 27523
rect 12265 27489 12299 27523
rect 13093 27489 13127 27523
rect 4813 27421 4847 27455
rect 6929 27421 6963 27455
rect 8493 27421 8527 27455
rect 9505 27421 9539 27455
rect 9597 27421 9631 27455
rect 9781 27421 9815 27455
rect 13277 27421 13311 27455
rect 15577 27421 15611 27455
rect 15669 27421 15703 27455
rect 15853 27421 15887 27455
rect 16681 27421 16715 27455
rect 16774 27421 16808 27455
rect 16957 27421 16991 27455
rect 17146 27421 17180 27455
rect 17405 27421 17439 27455
rect 17601 27421 17635 27455
rect 17693 27421 17727 27455
rect 17785 27421 17819 27455
rect 18153 27421 18187 27455
rect 18337 27421 18371 27455
rect 18429 27421 18463 27455
rect 18613 27421 18647 27455
rect 22937 27421 22971 27455
rect 23213 27421 23247 27455
rect 23489 27421 23523 27455
rect 23581 27421 23615 27455
rect 25513 27421 25547 27455
rect 25605 27421 25639 27455
rect 25789 27421 25823 27455
rect 27905 27421 27939 27455
rect 28181 27421 28215 27455
rect 29561 27421 29595 27455
rect 30021 27421 30055 27455
rect 30389 27421 30423 27455
rect 30482 27421 30516 27455
rect 30665 27421 30699 27455
rect 30895 27421 30929 27455
rect 33701 27421 33735 27455
rect 33977 27421 34011 27455
rect 10057 27353 10091 27387
rect 14473 27353 14507 27387
rect 17049 27353 17083 27387
rect 18061 27353 18095 27387
rect 18521 27353 18555 27387
rect 22753 27353 22787 27387
rect 23121 27353 23155 27387
rect 23397 27353 23431 27387
rect 26065 27353 26099 27387
rect 30757 27353 30791 27387
rect 6837 27285 6871 27319
rect 11529 27285 11563 27319
rect 11621 27285 11655 27319
rect 11989 27285 12023 27319
rect 14289 27285 14323 27319
rect 14381 27285 14415 27319
rect 17325 27285 17359 27319
rect 18797 27285 18831 27319
rect 27537 27285 27571 27319
rect 27813 27285 27847 27319
rect 27997 27285 28031 27319
rect 29653 27285 29687 27319
rect 29837 27285 29871 27319
rect 31033 27285 31067 27319
rect 33609 27285 33643 27319
rect 10241 27081 10275 27115
rect 16681 27081 16715 27115
rect 16957 27081 16991 27115
rect 18061 27081 18095 27115
rect 18797 27081 18831 27115
rect 22201 27081 22235 27115
rect 26985 27081 27019 27115
rect 12541 27013 12575 27047
rect 15485 27013 15519 27047
rect 22569 27013 22603 27047
rect 26341 27013 26375 27047
rect 29745 27013 29779 27047
rect 6653 26945 6687 26979
rect 10425 26945 10459 26979
rect 12265 26945 12299 26979
rect 12358 26945 12392 26979
rect 12633 26945 12667 26979
rect 12771 26945 12805 26979
rect 14473 26945 14507 26979
rect 14749 26945 14783 26979
rect 14933 26945 14967 26979
rect 15669 26945 15703 26979
rect 16865 26945 16899 26979
rect 17049 26945 17083 26979
rect 17693 26945 17727 26979
rect 17785 26945 17819 26979
rect 18981 26945 19015 26979
rect 19165 26945 19199 26979
rect 22385 26945 22419 26979
rect 22477 26945 22511 26979
rect 22753 26945 22787 26979
rect 26433 26945 26467 26979
rect 27169 26945 27203 26979
rect 27537 26945 27571 26979
rect 29469 26945 29503 26979
rect 31677 26945 31711 26979
rect 33149 26945 33183 26979
rect 33425 26945 33459 26979
rect 6929 26877 6963 26911
rect 8401 26877 8435 26911
rect 14657 26877 14691 26911
rect 26249 26877 26283 26911
rect 27813 26877 27847 26911
rect 33701 26877 33735 26911
rect 35449 26877 35483 26911
rect 14565 26809 14599 26843
rect 17233 26809 17267 26843
rect 26801 26809 26835 26843
rect 33333 26809 33367 26843
rect 12909 26741 12943 26775
rect 14289 26741 14323 26775
rect 17693 26741 17727 26775
rect 18981 26741 19015 26775
rect 29285 26741 29319 26775
rect 31217 26741 31251 26775
rect 31493 26741 31527 26775
rect 7757 26537 7791 26571
rect 13829 26537 13863 26571
rect 14473 26537 14507 26571
rect 17417 26537 17451 26571
rect 27813 26537 27847 26571
rect 30297 26537 30331 26571
rect 33241 26537 33275 26571
rect 15117 26469 15151 26503
rect 21373 26469 21407 26503
rect 25973 26469 26007 26503
rect 34897 26469 34931 26503
rect 7573 26401 7607 26435
rect 8677 26401 8711 26435
rect 28273 26401 28307 26435
rect 28365 26401 28399 26435
rect 29653 26401 29687 26435
rect 31309 26401 31343 26435
rect 33057 26401 33091 26435
rect 33885 26401 33919 26435
rect 35265 26401 35299 26435
rect 4537 26333 4571 26367
rect 4629 26333 4663 26367
rect 4813 26333 4847 26367
rect 7389 26333 7423 26367
rect 7941 26333 7975 26367
rect 8401 26333 8435 26367
rect 9137 26333 9171 26367
rect 13553 26333 13587 26367
rect 13645 26333 13679 26367
rect 13921 26333 13955 26367
rect 14657 26333 14691 26367
rect 15025 26333 15059 26367
rect 15301 26333 15335 26367
rect 15393 26333 15427 26367
rect 15669 26333 15703 26367
rect 16221 26333 16255 26367
rect 16865 26333 16899 26367
rect 17279 26333 17313 26367
rect 20821 26333 20855 26367
rect 21097 26333 21131 26367
rect 21189 26333 21223 26367
rect 23581 26333 23615 26367
rect 23857 26333 23891 26367
rect 25421 26333 25455 26367
rect 25605 26333 25639 26367
rect 25789 26333 25823 26367
rect 26249 26333 26283 26367
rect 26341 26333 26375 26367
rect 26525 26333 26559 26367
rect 26617 26333 26651 26367
rect 29837 26333 29871 26367
rect 30757 26333 30791 26367
rect 30849 26333 30883 26367
rect 31033 26333 31067 26367
rect 33609 26333 33643 26367
rect 34713 26333 34747 26367
rect 34989 26333 35023 26367
rect 5089 26265 5123 26299
rect 6837 26265 6871 26299
rect 8493 26265 8527 26299
rect 13369 26265 13403 26299
rect 14749 26265 14783 26299
rect 14841 26265 14875 26299
rect 15485 26265 15519 26299
rect 16037 26265 16071 26299
rect 16405 26265 16439 26299
rect 17049 26265 17083 26299
rect 17141 26265 17175 26299
rect 20269 26265 20303 26299
rect 20453 26265 20487 26299
rect 20637 26265 20671 26299
rect 21005 26265 21039 26299
rect 25697 26265 25731 26299
rect 28181 26265 28215 26299
rect 29929 26265 29963 26299
rect 33701 26265 33735 26299
rect 37013 26265 37047 26299
rect 6929 26197 6963 26231
rect 7297 26197 7331 26231
rect 8033 26197 8067 26231
rect 9045 26197 9079 26231
rect 23397 26197 23431 26231
rect 23765 26197 23799 26231
rect 26065 26197 26099 26231
rect 5457 25993 5491 26027
rect 16405 25993 16439 26027
rect 23949 25993 23983 26027
rect 25237 25993 25271 26027
rect 31585 25993 31619 26027
rect 32137 25993 32171 26027
rect 32597 25993 32631 26027
rect 34805 25993 34839 26027
rect 35265 25993 35299 26027
rect 19073 25925 19107 25959
rect 19533 25925 19567 25959
rect 20637 25925 20671 25959
rect 31953 25925 31987 25959
rect 1777 25857 1811 25891
rect 3065 25857 3099 25891
rect 5641 25857 5675 25891
rect 16221 25857 16255 25891
rect 18705 25857 18739 25891
rect 18797 25857 18831 25891
rect 18889 25857 18923 25891
rect 19324 25857 19358 25891
rect 19441 25857 19475 25891
rect 19688 25857 19722 25891
rect 19809 25857 19843 25891
rect 20453 25857 20487 25891
rect 20729 25857 20763 25891
rect 20821 25857 20855 25891
rect 22477 25857 22511 25891
rect 22661 25857 22695 25891
rect 22753 25857 22787 25891
rect 23121 25857 23155 25891
rect 23397 25857 23431 25891
rect 23857 25857 23891 25891
rect 24317 25857 24351 25891
rect 24593 25857 24627 25891
rect 24777 25857 24811 25891
rect 24869 25857 24903 25891
rect 24961 25857 24995 25891
rect 25513 25857 25547 25891
rect 25605 25857 25639 25891
rect 25697 25857 25731 25891
rect 25881 25857 25915 25891
rect 25973 25857 26007 25891
rect 26157 25857 26191 25891
rect 26249 25857 26283 25891
rect 26341 25857 26375 25891
rect 31493 25857 31527 25891
rect 31769 25857 31803 25891
rect 32505 25857 32539 25891
rect 32965 25857 32999 25891
rect 33149 25857 33183 25891
rect 33241 25857 33275 25891
rect 33333 25857 33367 25891
rect 34437 25857 34471 25891
rect 35081 25857 35115 25891
rect 35173 25857 35207 25891
rect 3341 25789 3375 25823
rect 3617 25789 3651 25823
rect 8677 25789 8711 25823
rect 8953 25789 8987 25823
rect 23765 25789 23799 25823
rect 24225 25789 24259 25823
rect 32689 25789 32723 25823
rect 34161 25789 34195 25823
rect 34345 25789 34379 25823
rect 18521 25721 18555 25755
rect 22569 25721 22603 25755
rect 23489 25721 23523 25755
rect 34989 25721 35023 25755
rect 1501 25653 1535 25687
rect 2881 25653 2915 25687
rect 5089 25653 5123 25687
rect 10425 25653 10459 25687
rect 19165 25653 19199 25687
rect 21005 25653 21039 25687
rect 22293 25653 22327 25687
rect 23673 25653 23707 25687
rect 24133 25653 24167 25687
rect 25329 25653 25363 25687
rect 26617 25653 26651 25687
rect 33609 25653 33643 25687
rect 3893 25449 3927 25483
rect 9045 25449 9079 25483
rect 22845 25449 22879 25483
rect 24777 25449 24811 25483
rect 11897 25381 11931 25415
rect 12817 25381 12851 25415
rect 16405 25381 16439 25415
rect 27813 25381 27847 25415
rect 2145 25313 2179 25347
rect 9873 25313 9907 25347
rect 12541 25313 12575 25347
rect 14841 25313 14875 25347
rect 17417 25313 17451 25347
rect 19073 25313 19107 25347
rect 21005 25313 21039 25347
rect 23489 25313 23523 25347
rect 1869 25245 1903 25279
rect 4077 25245 4111 25279
rect 7573 25245 7607 25279
rect 9229 25245 9263 25279
rect 9689 25245 9723 25279
rect 10149 25245 10183 25279
rect 12357 25245 12391 25279
rect 12955 25245 12989 25279
rect 13093 25245 13127 25279
rect 13313 25245 13347 25279
rect 13461 25245 13495 25279
rect 14565 25245 14599 25279
rect 15945 25245 15979 25279
rect 16680 25223 16714 25257
rect 16773 25245 16807 25279
rect 16865 25245 16899 25279
rect 17049 25245 17083 25279
rect 17233 25245 17267 25279
rect 18337 25245 18371 25279
rect 18521 25245 18555 25279
rect 18613 25245 18647 25279
rect 20729 25245 20763 25279
rect 20913 25245 20947 25279
rect 21235 25245 21269 25279
rect 21373 25245 21407 25279
rect 21465 25245 21499 25279
rect 21593 25245 21627 25279
rect 21741 25245 21775 25279
rect 22201 25245 22235 25279
rect 22349 25245 22383 25279
rect 22666 25245 22700 25279
rect 23029 25245 23063 25279
rect 24961 25245 24995 25279
rect 25053 25245 25087 25279
rect 25237 25245 25271 25279
rect 25329 25245 25363 25279
rect 27169 25245 27203 25279
rect 27262 25245 27296 25279
rect 27445 25245 27479 25279
rect 27634 25245 27668 25279
rect 28457 25245 28491 25279
rect 28733 25245 28767 25279
rect 29193 25245 29227 25279
rect 30021 25245 30055 25279
rect 30205 25245 30239 25279
rect 30297 25245 30331 25279
rect 30389 25245 30423 25279
rect 34345 25245 34379 25279
rect 34713 25245 34747 25279
rect 10425 25177 10459 25211
rect 12449 25177 12483 25211
rect 13185 25177 13219 25211
rect 22477 25177 22511 25211
rect 22569 25177 22603 25211
rect 27537 25177 27571 25211
rect 28549 25177 28583 25211
rect 28917 25177 28951 25211
rect 34989 25177 35023 25211
rect 36737 25177 36771 25211
rect 3617 25109 3651 25143
rect 7481 25109 7515 25143
rect 9321 25109 9355 25143
rect 9781 25109 9815 25143
rect 11989 25109 12023 25143
rect 16129 25109 16163 25143
rect 20545 25109 20579 25143
rect 21097 25109 21131 25143
rect 29101 25109 29135 25143
rect 30665 25109 30699 25143
rect 34529 25109 34563 25143
rect 4353 24905 4387 24939
rect 4721 24905 4755 24939
rect 9229 24905 9263 24939
rect 9597 24905 9631 24939
rect 10333 24905 10367 24939
rect 10609 24905 10643 24939
rect 12725 24905 12759 24939
rect 14289 24905 14323 24939
rect 18521 24905 18555 24939
rect 18705 24905 18739 24939
rect 21281 24905 21315 24939
rect 23397 24905 23431 24939
rect 27445 24905 27479 24939
rect 34253 24905 34287 24939
rect 12357 24837 12391 24871
rect 12817 24837 12851 24871
rect 13001 24837 13035 24871
rect 16221 24837 16255 24871
rect 18337 24837 18371 24871
rect 21097 24837 21131 24871
rect 21465 24837 21499 24871
rect 27353 24837 27387 24871
rect 30941 24837 30975 24871
rect 34621 24837 34655 24871
rect 5917 24769 5951 24803
rect 10425 24769 10459 24803
rect 10793 24769 10827 24803
rect 12173 24769 12207 24803
rect 12449 24769 12483 24803
rect 12541 24769 12575 24803
rect 14381 24769 14415 24803
rect 14841 24769 14875 24803
rect 15393 24769 15427 24803
rect 16681 24769 16715 24803
rect 16865 24769 16899 24803
rect 17233 24769 17267 24803
rect 21373 24769 21407 24803
rect 23489 24769 23523 24803
rect 24041 24769 24075 24803
rect 25881 24769 25915 24803
rect 26157 24769 26191 24803
rect 28641 24769 28675 24803
rect 28917 24769 28951 24803
rect 31125 24769 31159 24803
rect 31309 24769 31343 24803
rect 31585 24769 31619 24803
rect 31953 24769 31987 24803
rect 33057 24779 33091 24813
rect 33241 24769 33275 24803
rect 33517 24769 33551 24803
rect 1409 24701 1443 24735
rect 1685 24701 1719 24735
rect 4813 24701 4847 24735
rect 4997 24701 5031 24735
rect 7297 24701 7331 24735
rect 7573 24701 7607 24735
rect 9689 24701 9723 24735
rect 9873 24701 9907 24735
rect 15025 24701 15059 24735
rect 17325 24701 17359 24735
rect 17877 24701 17911 24735
rect 21649 24701 21683 24735
rect 24133 24701 24167 24735
rect 25789 24701 25823 24735
rect 27537 24701 27571 24735
rect 29193 24701 29227 24735
rect 33425 24701 33459 24735
rect 34713 24701 34747 24735
rect 34805 24701 34839 24735
rect 9045 24633 9079 24667
rect 26985 24633 27019 24667
rect 28825 24633 28859 24667
rect 3157 24565 3191 24599
rect 5733 24565 5767 24599
rect 13185 24565 13219 24599
rect 18521 24565 18555 24599
rect 25973 24565 26007 24599
rect 31217 24565 31251 24599
rect 33149 24565 33183 24599
rect 1777 24361 1811 24395
rect 3801 24361 3835 24395
rect 7941 24361 7975 24395
rect 13737 24361 13771 24395
rect 13921 24361 13955 24395
rect 18613 24361 18647 24395
rect 18797 24361 18831 24395
rect 27353 24361 27387 24395
rect 31769 24361 31803 24395
rect 15209 24293 15243 24327
rect 16865 24293 16899 24327
rect 18153 24293 18187 24327
rect 19901 24293 19935 24327
rect 20729 24293 20763 24327
rect 22109 24293 22143 24327
rect 33517 24293 33551 24327
rect 33701 24293 33735 24327
rect 34437 24293 34471 24327
rect 2973 24225 3007 24259
rect 4353 24225 4387 24259
rect 5273 24225 5307 24259
rect 5549 24225 5583 24259
rect 13001 24225 13035 24259
rect 16405 24225 16439 24259
rect 23305 24225 23339 24259
rect 25605 24225 25639 24259
rect 25881 24225 25915 24259
rect 28273 24225 28307 24259
rect 33057 24225 33091 24259
rect 1961 24157 1995 24191
rect 4169 24157 4203 24191
rect 8125 24157 8159 24191
rect 9137 24157 9171 24191
rect 12817 24157 12851 24191
rect 14289 24157 14323 24191
rect 14749 24157 14783 24191
rect 15209 24157 15243 24191
rect 15761 24157 15795 24191
rect 15945 24157 15979 24191
rect 16037 24157 16071 24191
rect 16163 24157 16197 24191
rect 17107 24157 17141 24191
rect 17233 24157 17267 24191
rect 17325 24157 17359 24191
rect 17509 24157 17543 24191
rect 17877 24157 17911 24191
rect 18153 24157 18187 24191
rect 18705 24157 18739 24191
rect 18935 24157 18969 24191
rect 19073 24157 19107 24191
rect 19533 24157 19567 24191
rect 19717 24157 19751 24191
rect 19993 24157 20027 24191
rect 20361 24157 20395 24191
rect 20453 24157 20487 24191
rect 20545 24157 20579 24191
rect 20821 24157 20855 24191
rect 22109 24157 22143 24191
rect 22937 24157 22971 24191
rect 23673 24157 23707 24191
rect 23949 24157 23983 24191
rect 24225 24157 24259 24191
rect 24777 24157 24811 24191
rect 25329 24157 25363 24191
rect 28181 24157 28215 24191
rect 28457 24157 28491 24191
rect 29561 24157 29595 24191
rect 29740 24157 29774 24191
rect 29837 24157 29871 24191
rect 29929 24157 29963 24191
rect 31401 24157 31435 24191
rect 31585 24157 31619 24191
rect 31677 24157 31711 24191
rect 32229 24157 32263 24191
rect 32413 24157 32447 24191
rect 32781 24157 32815 24191
rect 32873 24157 32907 24191
rect 33149 24157 33183 24191
rect 33241 24157 33275 24191
rect 33333 24157 33367 24191
rect 33609 24157 33643 24191
rect 33885 24157 33919 24191
rect 34069 24157 34103 24191
rect 34161 24157 34195 24191
rect 34345 24157 34379 24191
rect 2697 24089 2731 24123
rect 13553 24089 13587 24123
rect 20085 24089 20119 24123
rect 33517 24089 33551 24123
rect 33977 24089 34011 24123
rect 2329 24021 2363 24055
rect 2789 24021 2823 24055
rect 4261 24021 4295 24055
rect 7021 24021 7055 24055
rect 9045 24021 9079 24055
rect 12633 24021 12667 24055
rect 13763 24021 13797 24055
rect 18337 24021 18371 24055
rect 19257 24021 19291 24055
rect 19625 24021 19659 24055
rect 25237 24021 25271 24055
rect 30205 24021 30239 24055
rect 31493 24021 31527 24055
rect 32137 24021 32171 24055
rect 32413 24021 32447 24055
rect 32597 24021 32631 24055
rect 6377 23817 6411 23851
rect 6745 23817 6779 23851
rect 10425 23817 10459 23851
rect 14749 23817 14783 23851
rect 15761 23817 15795 23851
rect 18705 23817 18739 23851
rect 19349 23817 19383 23851
rect 19993 23817 20027 23851
rect 28641 23817 28675 23851
rect 29101 23817 29135 23851
rect 32229 23817 32263 23851
rect 13461 23749 13495 23783
rect 14289 23749 14323 23783
rect 14657 23749 14691 23783
rect 15025 23749 15059 23783
rect 16037 23749 16071 23783
rect 21097 23749 21131 23783
rect 22385 23749 22419 23783
rect 25881 23749 25915 23783
rect 27261 23749 27295 23783
rect 28733 23749 28767 23783
rect 5641 23681 5675 23715
rect 6837 23681 6871 23715
rect 8677 23681 8711 23715
rect 11161 23681 11195 23715
rect 12909 23681 12943 23715
rect 13001 23681 13035 23715
rect 14197 23681 14231 23715
rect 14841 23681 14875 23715
rect 15301 23681 15335 23715
rect 15485 23681 15519 23715
rect 15669 23681 15703 23715
rect 17325 23681 17359 23715
rect 17417 23681 17451 23715
rect 17969 23681 18003 23715
rect 18081 23681 18115 23715
rect 19073 23681 19107 23715
rect 19165 23681 19199 23715
rect 19441 23681 19475 23715
rect 19809 23681 19843 23715
rect 19901 23681 19935 23715
rect 20821 23681 20855 23715
rect 22569 23681 22603 23715
rect 23305 23681 23339 23715
rect 23673 23681 23707 23715
rect 23857 23681 23891 23715
rect 24685 23681 24719 23715
rect 25053 23681 25087 23715
rect 25145 23681 25179 23715
rect 26065 23681 26099 23715
rect 26157 23681 26191 23715
rect 27077 23681 27111 23715
rect 27353 23681 27387 23715
rect 27445 23681 27479 23715
rect 27721 23681 27755 23715
rect 27905 23681 27939 23715
rect 27997 23681 28031 23715
rect 28089 23681 28123 23715
rect 32137 23681 32171 23715
rect 33149 23681 33183 23715
rect 35541 23681 35575 23715
rect 6929 23613 6963 23647
rect 8953 23613 8987 23647
rect 15853 23613 15887 23647
rect 17233 23613 17267 23647
rect 17509 23613 17543 23647
rect 20269 23613 20303 23647
rect 22661 23613 22695 23647
rect 23213 23613 23247 23647
rect 28457 23613 28491 23647
rect 34989 23613 35023 23647
rect 35817 23613 35851 23647
rect 10609 23545 10643 23579
rect 18981 23545 19015 23579
rect 19533 23545 19567 23579
rect 20177 23545 20211 23579
rect 22201 23545 22235 23579
rect 24317 23545 24351 23579
rect 27629 23545 27663 23579
rect 28273 23545 28307 23579
rect 5549 23477 5583 23511
rect 12725 23477 12759 23511
rect 15117 23477 15151 23511
rect 15945 23477 15979 23511
rect 17693 23477 17727 23511
rect 17785 23477 17819 23511
rect 18245 23477 18279 23511
rect 33241 23477 33275 23511
rect 2237 23273 2271 23307
rect 2973 23273 3007 23307
rect 4261 23273 4295 23307
rect 4997 23273 5031 23307
rect 6285 23273 6319 23307
rect 6469 23273 6503 23307
rect 7021 23273 7055 23307
rect 8125 23273 8159 23307
rect 9321 23273 9355 23307
rect 14105 23273 14139 23307
rect 20453 23273 20487 23307
rect 20821 23273 20855 23307
rect 23857 23273 23891 23307
rect 34805 23273 34839 23307
rect 23489 23205 23523 23239
rect 5733 23137 5767 23171
rect 12817 23137 12851 23171
rect 15669 23137 15703 23171
rect 16221 23137 16255 23171
rect 18705 23137 18739 23171
rect 20545 23137 20579 23171
rect 22017 23137 22051 23171
rect 22753 23137 22787 23171
rect 35633 23137 35667 23171
rect 1961 23069 1995 23103
rect 2513 23069 2547 23103
rect 2605 23069 2639 23103
rect 2697 23069 2731 23103
rect 2881 23069 2915 23103
rect 3157 23069 3191 23103
rect 3341 23069 3375 23103
rect 3617 23069 3651 23103
rect 4445 23069 4479 23103
rect 4629 23069 4663 23103
rect 4905 23069 4939 23103
rect 5181 23069 5215 23103
rect 5641 23069 5675 23103
rect 5917 23069 5951 23103
rect 6193 23069 6227 23103
rect 6745 23069 6779 23103
rect 6929 23069 6963 23103
rect 7206 23047 7240 23081
rect 7665 23069 7699 23103
rect 7757 23069 7791 23103
rect 9505 23069 9539 23103
rect 9597 23069 9631 23103
rect 9873 23069 9907 23103
rect 10517 23069 10551 23103
rect 10609 23069 10643 23103
rect 10793 23069 10827 23103
rect 15209 23069 15243 23103
rect 15393 23069 15427 23103
rect 15761 23069 15795 23103
rect 16681 23069 16715 23103
rect 17049 23069 17083 23103
rect 17141 23069 17175 23103
rect 17417 23069 17451 23103
rect 17693 23069 17727 23103
rect 18245 23069 18279 23103
rect 18613 23069 18647 23103
rect 20453 23069 20487 23103
rect 21189 23069 21223 23103
rect 21741 23069 21775 23103
rect 22937 23069 22971 23103
rect 23397 23069 23431 23103
rect 23765 23069 23799 23103
rect 23949 23069 23983 23103
rect 24961 23069 24995 23103
rect 25237 23069 25271 23103
rect 25697 23069 25731 23103
rect 26065 23069 26099 23103
rect 29745 23069 29779 23103
rect 29929 23069 29963 23103
rect 32505 23069 32539 23103
rect 32781 23069 32815 23103
rect 32873 23069 32907 23103
rect 33057 23069 33091 23103
rect 34713 23069 34747 23103
rect 34989 23069 35023 23103
rect 35173 23069 35207 23103
rect 35265 23069 35299 23103
rect 35357 23069 35391 23103
rect 35725 23069 35759 23103
rect 35909 23069 35943 23103
rect 36185 23069 36219 23103
rect 36369 23069 36403 23103
rect 3249 23001 3283 23035
rect 3479 23001 3513 23035
rect 4537 23001 4571 23035
rect 4747 23001 4781 23035
rect 5273 23001 5307 23035
rect 5365 23001 5399 23035
rect 5483 23001 5517 23035
rect 6437 23001 6471 23035
rect 6653 23001 6687 23035
rect 7297 23001 7331 23035
rect 7389 23001 7423 23035
rect 7527 23001 7561 23035
rect 7941 23001 7975 23035
rect 9689 23001 9723 23035
rect 11069 23001 11103 23035
rect 14289 23001 14323 23035
rect 14473 23001 14507 23035
rect 14749 23001 14783 23035
rect 21005 23001 21039 23035
rect 25881 23001 25915 23035
rect 25973 23001 26007 23035
rect 30021 23001 30055 23035
rect 33241 23001 33275 23035
rect 1777 22933 1811 22967
rect 6101 22933 6135 22967
rect 6929 22933 6963 22967
rect 25421 22933 25455 22967
rect 26249 22933 26283 22967
rect 32321 22933 32355 22967
rect 32689 22933 32723 22967
rect 35541 22933 35575 22967
rect 36093 22933 36127 22967
rect 36277 22933 36311 22967
rect 2881 22729 2915 22763
rect 3433 22729 3467 22763
rect 3985 22729 4019 22763
rect 5089 22729 5123 22763
rect 5549 22729 5583 22763
rect 9505 22729 9539 22763
rect 11069 22729 11103 22763
rect 11529 22729 11563 22763
rect 11897 22729 11931 22763
rect 13001 22729 13035 22763
rect 13829 22729 13863 22763
rect 15301 22729 15335 22763
rect 15485 22729 15519 22763
rect 17969 22729 18003 22763
rect 20453 22729 20487 22763
rect 22109 22729 22143 22763
rect 24409 22729 24443 22763
rect 27537 22729 27571 22763
rect 27997 22729 28031 22763
rect 30297 22729 30331 22763
rect 32229 22729 32263 22763
rect 33701 22729 33735 22763
rect 37381 22729 37415 22763
rect 3617 22661 3651 22695
rect 5457 22661 5491 22695
rect 6561 22661 6595 22695
rect 8033 22661 8067 22695
rect 8217 22661 8251 22695
rect 13645 22661 13679 22695
rect 16129 22661 16163 22695
rect 16313 22661 16347 22695
rect 35173 22661 35207 22695
rect 36829 22661 36863 22695
rect 2789 22593 2823 22627
rect 2973 22593 3007 22627
rect 3801 22593 3835 22627
rect 3893 22593 3927 22627
rect 4077 22593 4111 22627
rect 5273 22593 5307 22627
rect 5549 22593 5583 22627
rect 5733 22593 5767 22627
rect 6377 22593 6411 22627
rect 7849 22593 7883 22627
rect 9689 22593 9723 22627
rect 9873 22593 9907 22627
rect 11253 22593 11287 22627
rect 12357 22593 12391 22627
rect 12541 22593 12575 22627
rect 12633 22593 12667 22627
rect 12725 22593 12759 22627
rect 13369 22593 13403 22627
rect 13553 22593 13587 22627
rect 14289 22593 14323 22627
rect 14657 22593 14691 22627
rect 15483 22593 15517 22627
rect 15945 22593 15979 22627
rect 17141 22593 17175 22627
rect 17325 22593 17359 22627
rect 17877 22593 17911 22627
rect 20729 22593 20763 22627
rect 22017 22593 22051 22627
rect 22201 22593 22235 22627
rect 22569 22593 22603 22627
rect 22661 22593 22695 22627
rect 23029 22593 23063 22627
rect 23397 22593 23431 22627
rect 23581 22593 23615 22627
rect 24041 22593 24075 22627
rect 24317 22593 24351 22627
rect 24501 22593 24535 22627
rect 25605 22593 25639 22627
rect 25789 22593 25823 22627
rect 26985 22593 27019 22627
rect 27169 22593 27203 22627
rect 27261 22593 27295 22627
rect 27353 22593 27387 22627
rect 27721 22593 27755 22627
rect 29653 22593 29687 22627
rect 29837 22593 29871 22627
rect 29929 22593 29963 22627
rect 30205 22593 30239 22627
rect 30389 22593 30423 22627
rect 30481 22593 30515 22627
rect 30665 22593 30699 22627
rect 32137 22593 32171 22627
rect 32321 22593 32355 22627
rect 32782 22593 32816 22627
rect 33149 22593 33183 22627
rect 33241 22593 33275 22627
rect 33425 22593 33459 22627
rect 33517 22593 33551 22627
rect 35357 22593 35391 22627
rect 35449 22593 35483 22627
rect 36093 22593 36127 22627
rect 36277 22593 36311 22627
rect 36369 22593 36403 22627
rect 36553 22593 36587 22627
rect 36645 22593 36679 22627
rect 37289 22593 37323 22627
rect 37657 22593 37691 22627
rect 6745 22525 6779 22559
rect 9965 22525 9999 22559
rect 11989 22525 12023 22559
rect 12173 22525 12207 22559
rect 16497 22525 16531 22559
rect 30021 22525 30055 22559
rect 32689 22525 32723 22559
rect 32873 22525 32907 22559
rect 32965 22525 32999 22559
rect 15853 22457 15887 22491
rect 23949 22457 23983 22491
rect 37841 22457 37875 22491
rect 25421 22389 25455 22423
rect 29469 22389 29503 22423
rect 30665 22389 30699 22423
rect 32505 22389 32539 22423
rect 35173 22389 35207 22423
rect 36093 22389 36127 22423
rect 36461 22389 36495 22423
rect 37013 22389 37047 22423
rect 3985 22185 4019 22219
rect 10333 22185 10367 22219
rect 12173 22185 12207 22219
rect 32873 22185 32907 22219
rect 4169 22117 4203 22151
rect 17049 22117 17083 22151
rect 19257 22117 19291 22151
rect 24225 22117 24259 22151
rect 27813 22117 27847 22151
rect 30757 22117 30791 22151
rect 32137 22117 32171 22151
rect 32505 22117 32539 22151
rect 10057 22049 10091 22083
rect 11621 22049 11655 22083
rect 12265 22049 12299 22083
rect 14473 22049 14507 22083
rect 16497 22049 16531 22083
rect 23673 22049 23707 22083
rect 25329 22049 25363 22083
rect 27261 22049 27295 22083
rect 30389 22049 30423 22083
rect 31309 22049 31343 22083
rect 32597 22049 32631 22083
rect 33149 22049 33183 22083
rect 33241 22049 33275 22083
rect 33333 22049 33367 22083
rect 35357 22049 35391 22083
rect 35725 22049 35759 22083
rect 35817 22049 35851 22083
rect 36001 22049 36035 22083
rect 37013 22049 37047 22083
rect 1961 21981 1995 22015
rect 4261 21981 4295 22015
rect 7757 21981 7791 22015
rect 10241 21981 10275 22015
rect 10425 21981 10459 22015
rect 12817 21981 12851 22015
rect 14841 21981 14875 22015
rect 15025 21981 15059 22015
rect 15485 21981 15519 22015
rect 15577 21981 15611 22015
rect 15853 21981 15887 22015
rect 16037 21981 16071 22015
rect 16405 21981 16439 22015
rect 16865 21981 16899 22015
rect 17049 21981 17083 22015
rect 17509 21981 17543 22015
rect 19441 21981 19475 22015
rect 19717 21981 19751 22015
rect 19993 21981 20027 22015
rect 20177 21981 20211 22015
rect 22201 21981 22235 22015
rect 22385 21981 22419 22015
rect 22753 21981 22787 22015
rect 22937 21981 22971 22015
rect 23581 21981 23615 22015
rect 24685 21981 24719 22015
rect 24869 21981 24903 22015
rect 24961 21981 24995 22015
rect 25053 21981 25087 22015
rect 25789 21981 25823 22015
rect 26209 21981 26243 22015
rect 27445 21981 27479 22015
rect 27721 21981 27755 22015
rect 27997 21981 28031 22015
rect 28365 21981 28399 22015
rect 28641 21981 28675 22015
rect 28825 21981 28859 22015
rect 28917 21981 28951 22015
rect 29009 21981 29043 22015
rect 31217 21981 31251 22015
rect 31861 21981 31895 22015
rect 31953 21981 31987 22015
rect 32137 21981 32171 22015
rect 32413 21981 32447 22015
rect 32689 21981 32723 22015
rect 33057 21981 33091 22015
rect 35081 21981 35115 22015
rect 35909 21981 35943 22015
rect 36829 21981 36863 22015
rect 3801 21913 3835 21947
rect 12449 21913 12483 21947
rect 22661 21913 22695 21947
rect 25973 21913 26007 21947
rect 26065 21913 26099 21947
rect 28181 21913 28215 21947
rect 28273 21913 28307 21947
rect 29837 21913 29871 21947
rect 31125 21913 31159 21947
rect 32229 21913 32263 21947
rect 35173 21913 35207 21947
rect 1777 21845 1811 21879
rect 4001 21845 4035 21879
rect 4353 21845 4387 21879
rect 8217 21845 8251 21879
rect 9413 21845 9447 21879
rect 9781 21845 9815 21879
rect 9873 21845 9907 21879
rect 11713 21845 11747 21879
rect 11805 21845 11839 21879
rect 12541 21845 12575 21879
rect 12633 21845 12667 21879
rect 16773 21845 16807 21879
rect 26358 21845 26392 21879
rect 27629 21845 27663 21879
rect 28549 21845 28583 21879
rect 29193 21845 29227 21879
rect 34713 21845 34747 21879
rect 35541 21845 35575 21879
rect 36645 21845 36679 21879
rect 3249 21641 3283 21675
rect 9137 21641 9171 21675
rect 9781 21641 9815 21675
rect 11529 21641 11563 21675
rect 11897 21641 11931 21675
rect 14933 21641 14967 21675
rect 17325 21641 17359 21675
rect 17693 21641 17727 21675
rect 18981 21641 19015 21675
rect 20177 21641 20211 21675
rect 22937 21641 22971 21675
rect 23581 21641 23615 21675
rect 27721 21641 27755 21675
rect 29929 21641 29963 21675
rect 32597 21641 32631 21675
rect 35265 21641 35299 21675
rect 35909 21641 35943 21675
rect 36461 21641 36495 21675
rect 1685 21573 1719 21607
rect 4563 21573 4597 21607
rect 5181 21573 5215 21607
rect 13829 21573 13863 21607
rect 23121 21573 23155 21607
rect 25053 21573 25087 21607
rect 25605 21573 25639 21607
rect 29745 21573 29779 21607
rect 33885 21573 33919 21607
rect 36369 21573 36403 21607
rect 3617 21505 3651 21539
rect 3709 21505 3743 21539
rect 4077 21505 4111 21539
rect 4261 21505 4295 21539
rect 4353 21505 4387 21539
rect 4445 21505 4479 21539
rect 4721 21505 4755 21539
rect 4997 21505 5031 21539
rect 5733 21505 5767 21539
rect 5825 21505 5859 21539
rect 5917 21505 5951 21539
rect 6101 21505 6135 21539
rect 9321 21505 9355 21539
rect 9413 21505 9447 21539
rect 9505 21505 9539 21539
rect 9689 21505 9723 21539
rect 9965 21505 9999 21539
rect 10057 21505 10091 21539
rect 10149 21505 10183 21539
rect 10333 21505 10367 21539
rect 13001 21505 13035 21539
rect 13277 21505 13311 21539
rect 13553 21505 13587 21539
rect 14289 21505 14323 21539
rect 14473 21505 14507 21539
rect 14565 21505 14599 21539
rect 15112 21505 15146 21539
rect 15209 21505 15243 21539
rect 15301 21505 15335 21539
rect 15484 21505 15518 21539
rect 15577 21505 15611 21539
rect 17509 21505 17543 21539
rect 17785 21505 17819 21539
rect 17877 21505 17911 21539
rect 19533 21505 19567 21539
rect 19901 21505 19935 21539
rect 20177 21505 20211 21539
rect 20361 21505 20395 21539
rect 23029 21505 23063 21539
rect 23397 21505 23431 21539
rect 24869 21505 24903 21539
rect 25145 21505 25179 21539
rect 25237 21505 25271 21539
rect 25697 21505 25731 21539
rect 27445 21505 27479 21539
rect 27629 21505 27663 21539
rect 27721 21505 27755 21539
rect 30021 21505 30055 21539
rect 30757 21505 30791 21539
rect 30941 21505 30975 21539
rect 32505 21505 32539 21539
rect 32689 21505 32723 21539
rect 33333 21505 33367 21539
rect 33425 21505 33459 21539
rect 33517 21505 33551 21539
rect 33701 21505 33735 21539
rect 33793 21505 33827 21539
rect 33977 21505 34011 21539
rect 35173 21505 35207 21539
rect 35817 21505 35851 21539
rect 36277 21505 36311 21539
rect 36737 21505 36771 21539
rect 1409 21437 1443 21471
rect 3157 21437 3191 21471
rect 3893 21437 3927 21471
rect 5365 21437 5399 21471
rect 6561 21437 6595 21471
rect 6837 21437 6871 21471
rect 11989 21437 12023 21471
rect 12173 21437 12207 21471
rect 13645 21437 13679 21471
rect 18061 21437 18095 21471
rect 18153 21437 18187 21471
rect 18521 21437 18555 21471
rect 19441 21437 19475 21471
rect 19809 21437 19843 21471
rect 23213 21437 23247 21471
rect 36001 21437 36035 21471
rect 8309 21369 8343 21403
rect 5457 21301 5491 21335
rect 23121 21301 23155 21335
rect 25421 21301 25455 21335
rect 29745 21301 29779 21335
rect 30941 21301 30975 21335
rect 33057 21301 33091 21335
rect 35449 21301 35483 21335
rect 4353 21097 4387 21131
rect 6929 21097 6963 21131
rect 9505 21097 9539 21131
rect 10149 21097 10183 21131
rect 14657 21097 14691 21131
rect 15485 21097 15519 21131
rect 16957 21097 16991 21131
rect 18429 21097 18463 21131
rect 18981 21097 19015 21131
rect 25053 21097 25087 21131
rect 26801 21097 26835 21131
rect 30573 21097 30607 21131
rect 7205 21029 7239 21063
rect 15209 21029 15243 21063
rect 21189 21029 21223 21063
rect 4077 20961 4111 20995
rect 4169 20961 4203 20995
rect 7665 20961 7699 20995
rect 7849 20961 7883 20995
rect 20269 20961 20303 20995
rect 25145 20961 25179 20995
rect 30665 20961 30699 20995
rect 1777 20893 1811 20927
rect 3893 20893 3927 20927
rect 3985 20893 4019 20927
rect 5457 20893 5491 20927
rect 7113 20893 7147 20927
rect 7573 20893 7607 20927
rect 8953 20893 8987 20927
rect 9321 20893 9355 20927
rect 9597 20893 9631 20927
rect 9965 20893 9999 20927
rect 14105 20893 14139 20927
rect 14381 20893 14415 20927
rect 14478 20893 14512 20927
rect 15393 20893 15427 20927
rect 15577 20893 15611 20927
rect 17136 20893 17170 20927
rect 17509 20893 17543 20927
rect 18554 20893 18588 20927
rect 19073 20893 19107 20927
rect 19349 20893 19383 20927
rect 19533 20893 19567 20927
rect 20177 20893 20211 20927
rect 20361 20893 20395 20927
rect 20545 20893 20579 20927
rect 20638 20893 20672 20927
rect 20821 20893 20855 20927
rect 21010 20893 21044 20927
rect 21373 20893 21407 20927
rect 21466 20893 21500 20927
rect 21838 20893 21872 20927
rect 22201 20893 22235 20927
rect 22385 20893 22419 20927
rect 22477 20893 22511 20927
rect 22569 20893 22603 20927
rect 25053 20893 25087 20927
rect 25329 20893 25363 20927
rect 26985 20893 27019 20927
rect 27077 20893 27111 20927
rect 27353 20893 27387 20927
rect 27629 20893 27663 20927
rect 27813 20893 27847 20927
rect 30389 20893 30423 20927
rect 34988 20903 35022 20937
rect 35081 20893 35115 20927
rect 35173 20893 35207 20927
rect 35357 20893 35391 20927
rect 35449 20893 35483 20927
rect 35633 20893 35667 20927
rect 37197 20893 37231 20927
rect 5273 20825 5307 20859
rect 5641 20825 5675 20859
rect 9137 20825 9171 20859
rect 9229 20825 9263 20859
rect 9781 20825 9815 20859
rect 9873 20825 9907 20859
rect 14289 20825 14323 20859
rect 14933 20825 14967 20859
rect 17233 20825 17267 20859
rect 17325 20825 17359 20859
rect 20913 20825 20947 20859
rect 21649 20825 21683 20859
rect 21741 20825 21775 20859
rect 27169 20825 27203 20859
rect 27445 20825 27479 20859
rect 34713 20825 34747 20859
rect 35541 20825 35575 20859
rect 37565 20825 37599 20859
rect 1501 20757 1535 20791
rect 18613 20757 18647 20791
rect 19441 20757 19475 20791
rect 22017 20757 22051 20791
rect 22845 20757 22879 20791
rect 24869 20757 24903 20791
rect 30205 20757 30239 20791
rect 37381 20757 37415 20791
rect 37841 20757 37875 20791
rect 3709 20553 3743 20587
rect 7573 20553 7607 20587
rect 14841 20553 14875 20587
rect 15669 20553 15703 20587
rect 18797 20553 18831 20587
rect 20177 20553 20211 20587
rect 21281 20553 21315 20587
rect 27813 20553 27847 20587
rect 35449 20553 35483 20587
rect 14657 20485 14691 20519
rect 19809 20485 19843 20519
rect 20545 20485 20579 20519
rect 27445 20485 27479 20519
rect 2789 20417 2823 20451
rect 3525 20417 3559 20451
rect 3801 20417 3835 20451
rect 7665 20417 7699 20451
rect 11713 20417 11747 20451
rect 15485 20417 15519 20451
rect 15577 20417 15611 20451
rect 18061 20417 18095 20451
rect 18153 20417 18187 20451
rect 18521 20417 18555 20451
rect 18613 20417 18647 20451
rect 19257 20417 19291 20451
rect 19993 20417 20027 20451
rect 20085 20417 20119 20451
rect 20361 20417 20395 20451
rect 20637 20417 20671 20451
rect 20730 20417 20764 20451
rect 20913 20417 20947 20451
rect 21005 20417 21039 20451
rect 21102 20417 21136 20451
rect 24317 20417 24351 20451
rect 24409 20417 24443 20451
rect 24593 20417 24627 20451
rect 25145 20417 25179 20451
rect 25789 20417 25823 20451
rect 25973 20417 26007 20451
rect 26065 20417 26099 20451
rect 26157 20417 26191 20451
rect 27261 20417 27295 20451
rect 27537 20417 27571 20451
rect 27629 20417 27663 20451
rect 28917 20417 28951 20451
rect 29101 20417 29135 20451
rect 29745 20417 29779 20451
rect 30297 20417 30331 20451
rect 30573 20417 30607 20451
rect 30757 20417 30791 20451
rect 31033 20417 31067 20451
rect 33149 20417 33183 20451
rect 35909 20417 35943 20451
rect 2881 20349 2915 20383
rect 3065 20349 3099 20383
rect 3341 20349 3375 20383
rect 7757 20349 7791 20383
rect 11621 20349 11655 20383
rect 14289 20349 14323 20383
rect 15945 20349 15979 20383
rect 17601 20349 17635 20383
rect 19165 20349 19199 20383
rect 24501 20349 24535 20383
rect 25329 20349 25363 20383
rect 29653 20349 29687 20383
rect 33241 20349 33275 20383
rect 35633 20349 35667 20383
rect 35725 20349 35759 20383
rect 35817 20349 35851 20383
rect 26341 20281 26375 20315
rect 30665 20281 30699 20315
rect 33517 20281 33551 20315
rect 2421 20213 2455 20247
rect 3893 20213 3927 20247
rect 7205 20213 7239 20247
rect 11989 20213 12023 20247
rect 14657 20213 14691 20247
rect 19441 20213 19475 20247
rect 19717 20213 19751 20247
rect 24133 20213 24167 20247
rect 24961 20213 24995 20247
rect 28917 20213 28951 20247
rect 30021 20213 30055 20247
rect 3801 20009 3835 20043
rect 9781 20009 9815 20043
rect 11621 20009 11655 20043
rect 13829 20009 13863 20043
rect 14749 20009 14783 20043
rect 15577 20009 15611 20043
rect 16405 20009 16439 20043
rect 16865 20009 16899 20043
rect 18889 20009 18923 20043
rect 20177 20009 20211 20043
rect 23121 20009 23155 20043
rect 23949 20009 23983 20043
rect 26341 20009 26375 20043
rect 26433 20009 26467 20043
rect 34897 20009 34931 20043
rect 36737 20009 36771 20043
rect 5089 19941 5123 19975
rect 8401 19941 8435 19975
rect 10425 19941 10459 19975
rect 12909 19941 12943 19975
rect 15853 19941 15887 19975
rect 16681 19941 16715 19975
rect 25605 19941 25639 19975
rect 29101 19941 29135 19975
rect 32321 19941 32355 19975
rect 35541 19941 35575 19975
rect 2973 19873 3007 19907
rect 4445 19873 4479 19907
rect 4813 19873 4847 19907
rect 5733 19873 5767 19907
rect 12173 19873 12207 19907
rect 19533 19873 19567 19907
rect 20269 19873 20303 19907
rect 23029 19873 23063 19907
rect 23857 19873 23891 19907
rect 24133 19873 24167 19907
rect 24869 19873 24903 19907
rect 25697 19873 25731 19907
rect 31033 19873 31067 19907
rect 31217 19873 31251 19907
rect 32045 19873 32079 19907
rect 36093 19873 36127 19907
rect 1961 19805 1995 19839
rect 3341 19805 3375 19839
rect 3985 19805 4019 19839
rect 4077 19805 4111 19839
rect 4721 19805 4755 19839
rect 5549 19805 5583 19839
rect 6193 19805 6227 19839
rect 6377 19805 6411 19839
rect 6561 19805 6595 19839
rect 6653 19805 6687 19839
rect 9229 19805 9263 19839
rect 9505 19805 9539 19839
rect 9597 19805 9631 19839
rect 9873 19805 9907 19839
rect 10149 19805 10183 19839
rect 10241 19805 10275 19839
rect 11989 19805 12023 19839
rect 12265 19805 12299 19839
rect 13185 19805 13219 19839
rect 13553 19805 13587 19839
rect 14105 19805 14139 19839
rect 14565 19805 14599 19839
rect 15209 19805 15243 19839
rect 15301 19805 15335 19839
rect 15669 19805 15703 19839
rect 16313 19805 16347 19839
rect 16405 19805 16439 19839
rect 16957 19805 16991 19839
rect 17417 19805 17451 19839
rect 17877 19805 17911 19839
rect 18153 19805 18187 19839
rect 18705 19805 18739 19839
rect 18973 19805 19007 19839
rect 19901 19805 19935 19839
rect 19993 19805 20027 19839
rect 20545 19805 20579 19839
rect 20637 19805 20671 19839
rect 20729 19805 20763 19839
rect 20913 19805 20947 19839
rect 23121 19805 23155 19839
rect 23673 19805 23707 19839
rect 24041 19805 24075 19839
rect 24225 19805 24259 19839
rect 24409 19805 24443 19839
rect 24593 19805 24627 19839
rect 24777 19805 24811 19839
rect 24961 19805 24995 19839
rect 25053 19805 25087 19839
rect 25421 19805 25455 19839
rect 26065 19805 26099 19839
rect 26157 19805 26191 19839
rect 26617 19805 26651 19839
rect 26709 19805 26743 19839
rect 26985 19805 27019 19839
rect 28457 19805 28491 19839
rect 28641 19805 28675 19839
rect 28917 19805 28951 19839
rect 29015 19805 29049 19839
rect 29193 19805 29227 19839
rect 29745 19805 29779 19839
rect 29837 19805 29871 19839
rect 30021 19805 30055 19839
rect 30113 19805 30147 19839
rect 30389 19805 30423 19839
rect 30665 19805 30699 19839
rect 31493 19805 31527 19839
rect 31953 19805 31987 19839
rect 33425 19805 33459 19839
rect 33609 19805 33643 19839
rect 35081 19805 35115 19839
rect 35173 19805 35207 19839
rect 35357 19805 35391 19839
rect 35449 19805 35483 19839
rect 36369 19805 36403 19839
rect 36553 19805 36587 19839
rect 36645 19805 36679 19839
rect 4169 19737 4203 19771
rect 4307 19737 4341 19771
rect 6285 19737 6319 19771
rect 6929 19737 6963 19771
rect 9413 19737 9447 19771
rect 10057 19737 10091 19771
rect 11621 19737 11655 19771
rect 13277 19737 13311 19771
rect 13645 19737 13679 19771
rect 19625 19737 19659 19771
rect 22845 19737 22879 19771
rect 23949 19737 23983 19771
rect 25237 19737 25271 19771
rect 25329 19737 25363 19771
rect 26801 19737 26835 19771
rect 28549 19737 28583 19771
rect 28825 19737 28859 19771
rect 36461 19737 36495 19771
rect 1777 19669 1811 19703
rect 5181 19669 5215 19703
rect 5641 19669 5675 19703
rect 6009 19669 6043 19703
rect 11437 19669 11471 19703
rect 12725 19669 12759 19703
rect 13461 19669 13495 19703
rect 23305 19669 23339 19703
rect 23489 19669 23523 19703
rect 24409 19669 24443 19703
rect 29561 19669 29595 19703
rect 33517 19669 33551 19703
rect 35909 19669 35943 19703
rect 36001 19669 36035 19703
rect 5917 19465 5951 19499
rect 7021 19465 7055 19499
rect 9321 19465 9355 19499
rect 12357 19465 12391 19499
rect 13185 19465 13219 19499
rect 19809 19465 19843 19499
rect 22661 19465 22695 19499
rect 23857 19465 23891 19499
rect 27813 19465 27847 19499
rect 30205 19465 30239 19499
rect 33793 19465 33827 19499
rect 33977 19465 34011 19499
rect 35909 19465 35943 19499
rect 1685 19397 1719 19431
rect 3893 19397 3927 19431
rect 8953 19397 8987 19431
rect 9045 19397 9079 19431
rect 13001 19397 13035 19431
rect 22201 19397 22235 19431
rect 23581 19397 23615 19431
rect 27445 19397 27479 19431
rect 27537 19397 27571 19431
rect 33333 19397 33367 19431
rect 1409 19329 1443 19363
rect 3525 19329 3559 19363
rect 3709 19329 3743 19363
rect 4169 19329 4203 19363
rect 7205 19329 7239 19363
rect 7941 19329 7975 19363
rect 8769 19329 8803 19363
rect 9137 19329 9171 19363
rect 9597 19329 9631 19363
rect 9781 19329 9815 19363
rect 11161 19329 11195 19363
rect 11345 19329 11379 19363
rect 11529 19329 11563 19363
rect 11897 19329 11931 19363
rect 11989 19329 12023 19363
rect 12265 19329 12299 19363
rect 12541 19329 12575 19363
rect 12633 19329 12667 19363
rect 13369 19329 13403 19363
rect 14289 19329 14323 19363
rect 14565 19329 14599 19363
rect 14749 19329 14783 19363
rect 16681 19329 16715 19363
rect 17141 19329 17175 19363
rect 17601 19329 17635 19363
rect 18153 19329 18187 19363
rect 19717 19329 19751 19363
rect 19901 19329 19935 19363
rect 22477 19329 22511 19363
rect 22753 19329 22787 19363
rect 24041 19329 24075 19363
rect 27281 19329 27315 19363
rect 27629 19329 27663 19363
rect 27905 19329 27939 19363
rect 28089 19329 28123 19363
rect 28273 19329 28307 19363
rect 29009 19329 29043 19363
rect 29193 19329 29227 19363
rect 29377 19329 29411 19363
rect 29469 19329 29503 19363
rect 29745 19329 29779 19363
rect 29837 19329 29871 19363
rect 30021 19329 30055 19363
rect 30205 19329 30239 19363
rect 32965 19329 32999 19363
rect 33149 19329 33183 19363
rect 33885 19329 33919 19363
rect 34161 19329 34195 19363
rect 34253 19329 34287 19363
rect 34437 19329 34471 19363
rect 34713 19329 34747 19363
rect 34897 19329 34931 19363
rect 35817 19329 35851 19363
rect 36001 19329 36035 19363
rect 4445 19261 4479 19295
rect 8309 19261 8343 19295
rect 9413 19261 9447 19295
rect 11805 19261 11839 19295
rect 13553 19261 13587 19295
rect 17969 19261 18003 19295
rect 22293 19261 22327 19295
rect 24317 19261 24351 19295
rect 29285 19261 29319 19295
rect 34805 19261 34839 19295
rect 3157 19193 3191 19227
rect 11713 19193 11747 19227
rect 14657 19193 14691 19227
rect 16773 19193 16807 19227
rect 33609 19193 33643 19227
rect 11345 19125 11379 19159
rect 12909 19125 12943 19159
rect 22477 19125 22511 19159
rect 24225 19125 24259 19159
rect 29653 19125 29687 19159
rect 33149 19125 33183 19159
rect 34621 19125 34655 19159
rect 4721 18921 4755 18955
rect 19809 18921 19843 18955
rect 20821 18921 20855 18955
rect 21005 18921 21039 18955
rect 22569 18921 22603 18955
rect 32965 18921 32999 18955
rect 17877 18853 17911 18887
rect 18337 18853 18371 18887
rect 22017 18853 22051 18887
rect 33609 18853 33643 18887
rect 3157 18785 3191 18819
rect 3341 18785 3375 18819
rect 5733 18785 5767 18819
rect 6101 18785 6135 18819
rect 10885 18785 10919 18819
rect 19349 18785 19383 18819
rect 19993 18785 20027 18819
rect 20177 18785 20211 18819
rect 20453 18785 20487 18819
rect 21833 18785 21867 18819
rect 22661 18785 22695 18819
rect 36737 18785 36771 18819
rect 4905 18717 4939 18751
rect 6009 18717 6043 18751
rect 10793 18717 10827 18751
rect 11805 18717 11839 18751
rect 11897 18717 11931 18751
rect 11989 18717 12023 18751
rect 12173 18717 12207 18751
rect 14381 18717 14415 18751
rect 14565 18717 14599 18751
rect 17693 18717 17727 18751
rect 17969 18717 18003 18751
rect 18061 18717 18095 18751
rect 18245 18717 18279 18751
rect 18521 18717 18555 18751
rect 18613 18717 18647 18751
rect 19257 18717 19291 18751
rect 19533 18717 19567 18751
rect 19625 18717 19659 18751
rect 20545 18717 20579 18751
rect 21557 18717 21591 18751
rect 21649 18717 21683 18751
rect 22385 18717 22419 18751
rect 31033 18717 31067 18751
rect 31217 18717 31251 18751
rect 31401 18717 31435 18751
rect 31585 18717 31619 18751
rect 32413 18717 32447 18751
rect 32505 18717 32539 18751
rect 32689 18717 32723 18751
rect 32781 18717 32815 18751
rect 33701 18717 33735 18751
rect 34989 18717 35023 18751
rect 36921 18717 36955 18751
rect 1409 18649 1443 18683
rect 1777 18649 1811 18683
rect 3065 18649 3099 18683
rect 5641 18649 5675 18683
rect 10701 18649 10735 18683
rect 11529 18649 11563 18683
rect 18337 18649 18371 18683
rect 21189 18649 21223 18683
rect 31493 18649 31527 18683
rect 34713 18649 34747 18683
rect 2697 18581 2731 18615
rect 6285 18581 6319 18615
rect 10333 18581 10367 18615
rect 14197 18581 14231 18615
rect 17509 18581 17543 18615
rect 18061 18581 18095 18615
rect 20989 18581 21023 18615
rect 22201 18581 22235 18615
rect 31217 18581 31251 18615
rect 34811 18581 34845 18615
rect 34897 18581 34931 18615
rect 37105 18581 37139 18615
rect 13921 18377 13955 18411
rect 15393 18377 15427 18411
rect 19441 18377 19475 18411
rect 25605 18377 25639 18411
rect 32781 18377 32815 18411
rect 34253 18377 34287 18411
rect 4353 18309 4387 18343
rect 9505 18309 9539 18343
rect 11253 18309 11287 18343
rect 12081 18309 12115 18343
rect 19901 18309 19935 18343
rect 32137 18309 32171 18343
rect 32965 18309 32999 18343
rect 33149 18309 33183 18343
rect 1869 18241 1903 18275
rect 2329 18241 2363 18275
rect 6193 18241 6227 18275
rect 11529 18241 11563 18275
rect 11713 18241 11747 18275
rect 12357 18241 12391 18275
rect 12541 18241 12575 18275
rect 14105 18241 14139 18275
rect 14289 18241 14323 18275
rect 14473 18241 14507 18275
rect 16957 18241 16991 18275
rect 17141 18241 17175 18275
rect 18797 18241 18831 18275
rect 18889 18241 18923 18275
rect 19257 18241 19291 18275
rect 19533 18241 19567 18275
rect 19626 18241 19660 18275
rect 22477 18241 22511 18275
rect 22753 18241 22787 18275
rect 23305 18241 23339 18275
rect 25053 18241 25087 18275
rect 25237 18241 25271 18275
rect 25329 18241 25363 18275
rect 25421 18241 25455 18275
rect 25881 18241 25915 18275
rect 27997 18241 28031 18275
rect 28181 18241 28215 18275
rect 29561 18241 29595 18275
rect 29745 18241 29779 18275
rect 30113 18241 30147 18275
rect 30665 18241 30699 18275
rect 31033 18241 31067 18275
rect 31217 18241 31251 18275
rect 31401 18241 31435 18275
rect 31493 18241 31527 18275
rect 31677 18241 31711 18275
rect 31861 18241 31895 18275
rect 32873 18241 32907 18275
rect 34345 18241 34379 18275
rect 34805 18241 34839 18275
rect 34989 18241 35023 18275
rect 35173 18241 35207 18275
rect 36921 18241 36955 18275
rect 37565 18241 37599 18275
rect 1685 18173 1719 18207
rect 2145 18173 2179 18207
rect 5917 18173 5951 18207
rect 7573 18173 7607 18207
rect 7849 18173 7883 18207
rect 12173 18173 12207 18207
rect 14749 18173 14783 18207
rect 15577 18173 15611 18207
rect 15669 18173 15703 18207
rect 16037 18173 16071 18207
rect 22937 18173 22971 18207
rect 25789 18173 25823 18207
rect 30481 18173 30515 18207
rect 32505 18173 32539 18207
rect 32597 18173 32631 18207
rect 34069 18173 34103 18207
rect 11713 18105 11747 18139
rect 23581 18105 23615 18139
rect 26249 18105 26283 18139
rect 33149 18105 33183 18139
rect 34713 18105 34747 18139
rect 2053 18037 2087 18071
rect 2513 18037 2547 18071
rect 3065 18037 3099 18071
rect 9321 18037 9355 18071
rect 18429 18037 18463 18071
rect 19165 18037 19199 18071
rect 28089 18037 28123 18071
rect 29561 18037 29595 18071
rect 34897 18037 34931 18071
rect 37105 18037 37139 18071
rect 37841 18037 37875 18071
rect 2053 17833 2087 17867
rect 2973 17833 3007 17867
rect 7849 17833 7883 17867
rect 8033 17833 8067 17867
rect 11345 17833 11379 17867
rect 12449 17833 12483 17867
rect 12817 17833 12851 17867
rect 15301 17833 15335 17867
rect 20637 17833 20671 17867
rect 22937 17833 22971 17867
rect 27353 17833 27387 17867
rect 31309 17833 31343 17867
rect 32137 17833 32171 17867
rect 8953 17765 8987 17799
rect 11253 17765 11287 17799
rect 16037 17765 16071 17799
rect 23949 17765 23983 17799
rect 25605 17765 25639 17799
rect 26617 17765 26651 17799
rect 34069 17765 34103 17799
rect 1593 17697 1627 17731
rect 3985 17697 4019 17731
rect 9413 17697 9447 17731
rect 9505 17697 9539 17731
rect 10057 17697 10091 17731
rect 10885 17697 10919 17731
rect 11805 17697 11839 17731
rect 11989 17697 12023 17731
rect 12541 17697 12575 17731
rect 14657 17697 14691 17731
rect 15485 17697 15519 17731
rect 23489 17697 23523 17731
rect 24685 17697 24719 17731
rect 24961 17697 24995 17731
rect 25145 17697 25179 17731
rect 26341 17697 26375 17731
rect 26985 17697 27019 17731
rect 27721 17697 27755 17731
rect 1777 17629 1811 17663
rect 2237 17629 2271 17663
rect 3249 17629 3283 17663
rect 3341 17629 3375 17663
rect 3433 17629 3467 17663
rect 3617 17629 3651 17663
rect 6101 17629 6135 17663
rect 8217 17629 8251 17663
rect 10149 17629 10183 17663
rect 10425 17629 10459 17663
rect 11069 17629 11103 17663
rect 11253 17629 11287 17663
rect 12633 17629 12667 17663
rect 12725 17629 12759 17663
rect 12909 17629 12943 17663
rect 13009 17629 13043 17663
rect 13185 17629 13219 17663
rect 13737 17629 13771 17663
rect 13921 17629 13955 17663
rect 14289 17629 14323 17663
rect 15577 17629 15611 17663
rect 15853 17629 15887 17663
rect 16267 17629 16301 17663
rect 16405 17629 16439 17663
rect 16497 17629 16531 17663
rect 16681 17629 16715 17663
rect 17417 17629 17451 17663
rect 17693 17629 17727 17663
rect 17877 17629 17911 17663
rect 18061 17629 18095 17663
rect 18153 17629 18187 17663
rect 18245 17629 18279 17663
rect 18429 17629 18463 17663
rect 18797 17629 18831 17663
rect 18981 17629 19015 17663
rect 20361 17629 20395 17663
rect 22293 17629 22327 17663
rect 22477 17629 22511 17663
rect 22569 17629 22603 17663
rect 22661 17629 22695 17663
rect 23581 17629 23615 17663
rect 24593 17629 24627 17663
rect 25237 17629 25271 17663
rect 26249 17629 26283 17663
rect 27077 17629 27111 17663
rect 27905 17629 27939 17663
rect 28365 17629 28399 17663
rect 28549 17629 28583 17663
rect 29193 17629 29227 17663
rect 29561 17629 29595 17663
rect 29745 17629 29779 17663
rect 29837 17629 29871 17663
rect 29929 17629 29963 17663
rect 30297 17629 30331 17663
rect 30481 17629 30515 17663
rect 31217 17629 31251 17663
rect 32045 17629 32079 17663
rect 33793 17629 33827 17663
rect 34069 17629 34103 17663
rect 4261 17561 4295 17595
rect 6377 17561 6411 17595
rect 11713 17561 11747 17595
rect 15945 17561 15979 17595
rect 20545 17561 20579 17595
rect 1961 17493 1995 17527
rect 5733 17493 5767 17527
rect 9321 17493 9355 17527
rect 12265 17493 12299 17527
rect 13001 17493 13035 17527
rect 13645 17493 13679 17527
rect 17509 17493 17543 17527
rect 18613 17493 18647 17527
rect 18889 17493 18923 17527
rect 30205 17493 30239 17527
rect 30389 17493 30423 17527
rect 33885 17493 33919 17527
rect 3433 17289 3467 17323
rect 4261 17289 4295 17323
rect 4537 17289 4571 17323
rect 6561 17289 6595 17323
rect 6929 17289 6963 17323
rect 7389 17289 7423 17323
rect 11989 17289 12023 17323
rect 14013 17289 14047 17323
rect 28365 17289 28399 17323
rect 29193 17289 29227 17323
rect 33149 17289 33183 17323
rect 33993 17289 34027 17323
rect 34161 17289 34195 17323
rect 4905 17221 4939 17255
rect 5917 17221 5951 17255
rect 9965 17221 9999 17255
rect 19901 17221 19935 17255
rect 19993 17221 20027 17255
rect 20361 17221 20395 17255
rect 28273 17221 28307 17255
rect 28533 17221 28567 17255
rect 28733 17221 28767 17255
rect 31677 17221 31711 17255
rect 33793 17221 33827 17255
rect 3065 17153 3099 17187
rect 3249 17153 3283 17187
rect 4445 17153 4479 17187
rect 5733 17153 5767 17187
rect 6745 17153 6779 17187
rect 7297 17153 7331 17187
rect 8953 17153 8987 17187
rect 9137 17153 9171 17187
rect 10240 17175 10274 17209
rect 10332 17175 10366 17209
rect 10425 17153 10459 17187
rect 10609 17153 10643 17187
rect 11989 17153 12023 17187
rect 12173 17153 12207 17187
rect 12265 17153 12299 17187
rect 12449 17153 12483 17187
rect 16681 17153 16715 17187
rect 16865 17153 16899 17187
rect 19625 17153 19659 17187
rect 19718 17153 19752 17187
rect 20090 17153 20124 17187
rect 20637 17153 20671 17187
rect 20729 17153 20763 17187
rect 20826 17153 20860 17187
rect 21005 17153 21039 17187
rect 22385 17153 22419 17187
rect 22937 17153 22971 17187
rect 23489 17153 23523 17187
rect 27997 17153 28031 17187
rect 28089 17153 28123 17187
rect 29009 17153 29043 17187
rect 29193 17153 29227 17187
rect 29561 17153 29595 17187
rect 31861 17153 31895 17187
rect 31953 17153 31987 17187
rect 32412 17153 32446 17187
rect 32873 17153 32907 17187
rect 33057 17153 33091 17187
rect 34437 17153 34471 17187
rect 34897 17153 34931 17187
rect 4997 17085 5031 17119
rect 5089 17085 5123 17119
rect 7481 17085 7515 17119
rect 12357 17085 12391 17119
rect 14473 17085 14507 17119
rect 22477 17085 22511 17119
rect 22753 17085 22787 17119
rect 32321 17085 32355 17119
rect 32505 17085 32539 17119
rect 32597 17085 32631 17119
rect 32781 17085 32815 17119
rect 34529 17085 34563 17119
rect 34989 17085 35023 17119
rect 35173 17085 35207 17119
rect 14197 17017 14231 17051
rect 28273 17017 28307 17051
rect 31677 17017 31711 17051
rect 6101 16949 6135 16983
rect 9321 16949 9355 16983
rect 16681 16949 16715 16983
rect 17049 16949 17083 16983
rect 20269 16949 20303 16983
rect 28549 16949 28583 16983
rect 33977 16949 34011 16983
rect 34437 16949 34471 16983
rect 34805 16949 34839 16983
rect 35081 16949 35115 16983
rect 16497 16745 16531 16779
rect 16681 16745 16715 16779
rect 30113 16745 30147 16779
rect 31217 16745 31251 16779
rect 32137 16745 32171 16779
rect 35173 16745 35207 16779
rect 35449 16745 35483 16779
rect 3801 16677 3835 16711
rect 8401 16677 8435 16711
rect 34345 16677 34379 16711
rect 34437 16677 34471 16711
rect 35357 16677 35391 16711
rect 2789 16609 2823 16643
rect 2973 16609 3007 16643
rect 4445 16609 4479 16643
rect 9137 16609 9171 16643
rect 16129 16609 16163 16643
rect 23213 16609 23247 16643
rect 23505 16609 23539 16643
rect 23949 16609 23983 16643
rect 25605 16609 25639 16643
rect 34253 16609 34287 16643
rect 35541 16609 35575 16643
rect 1961 16541 1995 16575
rect 2237 16541 2271 16575
rect 3985 16541 4019 16575
rect 4169 16541 4203 16575
rect 4529 16541 4563 16575
rect 8585 16541 8619 16575
rect 8769 16541 8803 16575
rect 14749 16541 14783 16575
rect 15393 16541 15427 16575
rect 16957 16541 16991 16575
rect 17233 16541 17267 16575
rect 17601 16541 17635 16575
rect 17969 16541 18003 16575
rect 18245 16541 18279 16575
rect 18337 16541 18371 16575
rect 18613 16541 18647 16575
rect 20269 16541 20303 16575
rect 20362 16541 20396 16575
rect 20637 16541 20671 16575
rect 20775 16541 20809 16575
rect 21005 16541 21039 16575
rect 21373 16541 21407 16575
rect 21833 16541 21867 16575
rect 22293 16541 22327 16575
rect 25237 16541 25271 16575
rect 25421 16541 25455 16575
rect 26065 16541 26099 16575
rect 30021 16541 30055 16575
rect 30205 16541 30239 16575
rect 30573 16541 30607 16575
rect 30757 16541 30791 16575
rect 31401 16541 31435 16575
rect 32321 16541 32355 16575
rect 34528 16519 34562 16553
rect 35449 16541 35483 16575
rect 4077 16473 4111 16507
rect 4307 16473 4341 16507
rect 9413 16473 9447 16507
rect 16773 16473 16807 16507
rect 19073 16473 19107 16507
rect 20545 16473 20579 16507
rect 22109 16473 22143 16507
rect 22845 16473 22879 16507
rect 23305 16473 23339 16507
rect 23765 16473 23799 16507
rect 26249 16473 26283 16507
rect 32505 16473 32539 16507
rect 34989 16473 35023 16507
rect 1777 16405 1811 16439
rect 2053 16405 2087 16439
rect 2329 16405 2363 16439
rect 2697 16405 2731 16439
rect 4629 16405 4663 16439
rect 10885 16405 10919 16439
rect 16497 16405 16531 16439
rect 17141 16405 17175 16439
rect 20913 16405 20947 16439
rect 23397 16405 23431 16439
rect 26433 16405 26467 16439
rect 30757 16405 30791 16439
rect 35189 16405 35223 16439
rect 35817 16405 35851 16439
rect 3893 16201 3927 16235
rect 4061 16201 4095 16235
rect 5181 16201 5215 16235
rect 9505 16201 9539 16235
rect 9781 16201 9815 16235
rect 10149 16201 10183 16235
rect 14473 16201 14507 16235
rect 16865 16201 16899 16235
rect 17709 16201 17743 16235
rect 17877 16201 17911 16235
rect 20729 16201 20763 16235
rect 21465 16201 21499 16235
rect 29285 16201 29319 16235
rect 30481 16201 30515 16235
rect 30849 16201 30883 16235
rect 34989 16201 35023 16235
rect 1685 16133 1719 16167
rect 4261 16133 4295 16167
rect 10241 16133 10275 16167
rect 17509 16133 17543 16167
rect 18797 16133 18831 16167
rect 20361 16133 20395 16167
rect 20561 16133 20595 16167
rect 23029 16133 23063 16167
rect 29395 16133 29429 16167
rect 29561 16133 29595 16167
rect 31033 16133 31067 16167
rect 31217 16133 31251 16167
rect 5549 16065 5583 16099
rect 9689 16065 9723 16099
rect 12265 16065 12299 16099
rect 12357 16065 12391 16099
rect 14013 16065 14047 16099
rect 14289 16065 14323 16099
rect 16957 16065 16991 16099
rect 17049 16065 17083 16099
rect 17969 16065 18003 16099
rect 18153 16065 18187 16099
rect 18245 16065 18279 16099
rect 18337 16065 18371 16099
rect 20269 16065 20303 16099
rect 21281 16065 21315 16099
rect 22845 16065 22879 16099
rect 23121 16065 23155 16099
rect 23213 16065 23247 16099
rect 24685 16065 24719 16099
rect 25237 16065 25271 16099
rect 26249 16065 26283 16099
rect 26341 16065 26375 16099
rect 27077 16065 27111 16099
rect 27353 16065 27387 16099
rect 29101 16065 29135 16099
rect 29276 16065 29310 16099
rect 30113 16065 30147 16099
rect 30665 16065 30699 16099
rect 30941 16065 30975 16099
rect 34897 16065 34931 16099
rect 35173 16065 35207 16099
rect 37657 16065 37691 16099
rect 1409 15997 1443 16031
rect 5641 15997 5675 16031
rect 5825 15997 5859 16031
rect 10333 15997 10367 16031
rect 12541 15997 12575 16031
rect 21005 15997 21039 16031
rect 26525 15997 26559 16031
rect 27261 15997 27295 16031
rect 29745 15997 29779 16031
rect 29929 15997 29963 16031
rect 11897 15929 11931 15963
rect 14105 15929 14139 15963
rect 17233 15929 17267 15963
rect 27169 15929 27203 15963
rect 3157 15861 3191 15895
rect 4077 15861 4111 15895
rect 16681 15861 16715 15895
rect 17693 15861 17727 15895
rect 18613 15861 18647 15895
rect 18889 15861 18923 15895
rect 20177 15861 20211 15895
rect 20545 15861 20579 15895
rect 21097 15861 21131 15895
rect 23397 15861 23431 15895
rect 25697 15861 25731 15895
rect 27537 15861 27571 15895
rect 30297 15861 30331 15895
rect 31401 15861 31435 15895
rect 35173 15861 35207 15895
rect 37841 15861 37875 15895
rect 1501 15657 1535 15691
rect 3801 15657 3835 15691
rect 4997 15657 5031 15691
rect 7941 15657 7975 15691
rect 10241 15657 10275 15691
rect 14289 15657 14323 15691
rect 14749 15657 14783 15691
rect 18153 15657 18187 15691
rect 26341 15657 26375 15691
rect 32321 15657 32355 15691
rect 32781 15657 32815 15691
rect 33241 15657 33275 15691
rect 35173 15657 35207 15691
rect 35449 15657 35483 15691
rect 26617 15589 26651 15623
rect 32413 15589 32447 15623
rect 4077 15521 4111 15555
rect 4537 15521 4571 15555
rect 6193 15521 6227 15555
rect 11529 15521 11563 15555
rect 15485 15521 15519 15555
rect 15761 15521 15795 15555
rect 15853 15521 15887 15555
rect 18797 15521 18831 15555
rect 20821 15521 20855 15555
rect 27721 15521 27755 15555
rect 27997 15521 28031 15555
rect 31861 15521 31895 15555
rect 32229 15521 32263 15555
rect 33333 15521 33367 15555
rect 34805 15521 34839 15555
rect 35633 15521 35667 15555
rect 1777 15453 1811 15487
rect 3985 15453 4019 15487
rect 4169 15453 4203 15487
rect 4261 15453 4295 15487
rect 4629 15453 4663 15487
rect 8953 15453 8987 15487
rect 11345 15453 11379 15487
rect 11897 15453 11931 15487
rect 14197 15453 14231 15487
rect 14565 15453 14599 15487
rect 15669 15453 15703 15487
rect 15945 15453 15979 15487
rect 16121 15455 16155 15489
rect 16313 15453 16347 15487
rect 18981 15453 19015 15487
rect 19073 15453 19107 15487
rect 19349 15453 19383 15487
rect 19993 15453 20027 15487
rect 20729 15453 20763 15487
rect 22937 15453 22971 15487
rect 23121 15453 23155 15487
rect 23397 15453 23431 15487
rect 23673 15453 23707 15487
rect 23765 15453 23799 15487
rect 24501 15453 24535 15487
rect 24777 15453 24811 15487
rect 24961 15453 24995 15487
rect 25237 15453 25271 15487
rect 25421 15453 25455 15487
rect 25973 15453 26007 15487
rect 26157 15453 26191 15487
rect 26433 15453 26467 15487
rect 27629 15453 27663 15487
rect 28181 15453 28215 15487
rect 28457 15453 28491 15487
rect 28641 15453 28675 15487
rect 28733 15453 28767 15487
rect 29653 15453 29687 15487
rect 29837 15453 29871 15487
rect 31493 15453 31527 15487
rect 31677 15453 31711 15487
rect 32505 15453 32539 15487
rect 33425 15453 33459 15487
rect 34897 15453 34931 15487
rect 35725 15453 35759 15487
rect 6469 15385 6503 15419
rect 12173 15385 12207 15419
rect 13921 15385 13955 15419
rect 18245 15385 18279 15419
rect 18429 15385 18463 15419
rect 32749 15385 32783 15419
rect 32965 15385 32999 15419
rect 10977 15317 11011 15351
rect 11437 15317 11471 15351
rect 16129 15317 16163 15351
rect 18613 15317 18647 15351
rect 19349 15317 19383 15351
rect 25605 15317 25639 15351
rect 27261 15317 27295 15351
rect 28365 15317 28399 15351
rect 30665 15317 30699 15351
rect 32597 15317 32631 15351
rect 33057 15317 33091 15351
rect 2973 15113 3007 15147
rect 3709 15113 3743 15147
rect 4077 15113 4111 15147
rect 6653 15113 6687 15147
rect 7573 15113 7607 15147
rect 11989 15113 12023 15147
rect 13921 15113 13955 15147
rect 15761 15113 15795 15147
rect 27077 15113 27111 15147
rect 34345 15113 34379 15147
rect 4905 15045 4939 15079
rect 9045 15045 9079 15079
rect 11897 15045 11931 15079
rect 14749 15045 14783 15079
rect 15025 15045 15059 15079
rect 29009 15045 29043 15079
rect 2881 14977 2915 15011
rect 3433 14977 3467 15011
rect 3617 14977 3651 15011
rect 4721 14977 4755 15011
rect 6837 14977 6871 15011
rect 7481 14977 7515 15011
rect 8125 14977 8159 15011
rect 8401 14977 8435 15011
rect 10517 14977 10551 15011
rect 13001 14977 13035 15011
rect 13369 14977 13403 15011
rect 14105 14977 14139 15011
rect 14197 14977 14231 15011
rect 14289 14977 14323 15011
rect 14473 14977 14507 15011
rect 14565 14977 14599 15011
rect 14841 14977 14875 15011
rect 15117 14977 15151 15011
rect 15485 14977 15519 15011
rect 15577 14977 15611 15011
rect 16221 14977 16255 15011
rect 16497 14977 16531 15011
rect 16865 14977 16899 15011
rect 17049 14977 17083 15011
rect 17141 14977 17175 15011
rect 17417 14977 17451 15011
rect 17693 14977 17727 15011
rect 18797 14977 18831 15011
rect 19165 14977 19199 15011
rect 19533 14977 19567 15011
rect 20085 14977 20119 15011
rect 20177 14977 20211 15011
rect 20361 14977 20395 15011
rect 22017 14977 22051 15011
rect 22201 14977 22235 15011
rect 22661 14977 22695 15011
rect 23213 14977 23247 15011
rect 25513 14977 25547 15011
rect 25697 14977 25731 15011
rect 25789 14977 25823 15011
rect 25973 14977 26007 15011
rect 26985 14977 27019 15011
rect 27261 14977 27295 15011
rect 27813 14977 27847 15011
rect 28089 14977 28123 15011
rect 28273 14977 28307 15011
rect 28457 14977 28491 15011
rect 28549 14977 28583 15011
rect 28641 14977 28675 15011
rect 28825 14977 28859 15011
rect 30665 14977 30699 15011
rect 30849 14977 30883 15011
rect 30941 14977 30975 15011
rect 31125 14977 31159 15011
rect 33057 14977 33091 15011
rect 33977 14977 34011 15011
rect 3157 14909 3191 14943
rect 4169 14909 4203 14943
rect 4261 14909 4295 14943
rect 4537 14909 4571 14943
rect 7665 14909 7699 14943
rect 7941 14909 7975 14943
rect 8309 14909 8343 14943
rect 9505 14909 9539 14943
rect 9597 14909 9631 14943
rect 12173 14909 12207 14943
rect 18153 14909 18187 14943
rect 21833 14909 21867 14943
rect 27909 14909 27943 14943
rect 32965 14909 32999 14943
rect 33885 14909 33919 14943
rect 7113 14841 7147 14875
rect 9045 14841 9079 14875
rect 11529 14841 11563 14875
rect 14841 14841 14875 14875
rect 15945 14841 15979 14875
rect 18797 14841 18831 14875
rect 27445 14841 27479 14875
rect 27997 14841 28031 14875
rect 30849 14841 30883 14875
rect 33425 14841 33459 14875
rect 2513 14773 2547 14807
rect 3617 14773 3651 14807
rect 8677 14773 8711 14807
rect 8861 14773 8895 14807
rect 9781 14773 9815 14807
rect 10333 14773 10367 14807
rect 12541 14773 12575 14807
rect 16405 14773 16439 14807
rect 20545 14773 20579 14807
rect 25605 14773 25639 14807
rect 25973 14773 26007 14807
rect 27629 14773 27663 14807
rect 31033 14773 31067 14807
rect 3157 14569 3191 14603
rect 4077 14569 4111 14603
rect 7389 14569 7423 14603
rect 13461 14569 13495 14603
rect 16589 14569 16623 14603
rect 17049 14569 17083 14603
rect 17417 14569 17451 14603
rect 19625 14569 19659 14603
rect 22293 14569 22327 14603
rect 23765 14569 23799 14603
rect 31953 14569 31987 14603
rect 10149 14433 10183 14467
rect 11897 14433 11931 14467
rect 12817 14433 12851 14467
rect 13001 14433 13035 14467
rect 15577 14433 15611 14467
rect 18061 14433 18095 14467
rect 21005 14433 21039 14467
rect 21649 14433 21683 14467
rect 23305 14433 23339 14467
rect 23397 14433 23431 14467
rect 30205 14433 30239 14467
rect 1409 14365 1443 14399
rect 4077 14365 4111 14399
rect 4261 14365 4295 14399
rect 5641 14365 5675 14399
rect 8953 14365 8987 14399
rect 9137 14365 9171 14399
rect 9229 14365 9263 14399
rect 9321 14365 9355 14399
rect 9873 14365 9907 14399
rect 15301 14365 15335 14399
rect 16589 14365 16623 14399
rect 16773 14365 16807 14399
rect 17049 14365 17083 14399
rect 17227 14365 17261 14399
rect 17325 14365 17359 14399
rect 17969 14365 18003 14399
rect 18153 14365 18187 14399
rect 19901 14365 19935 14399
rect 20269 14365 20303 14399
rect 20545 14365 20579 14399
rect 21281 14365 21315 14399
rect 22017 14365 22051 14399
rect 22661 14365 22695 14399
rect 23581 14365 23615 14399
rect 30389 14365 30423 14399
rect 31217 14365 31251 14399
rect 31401 14365 31435 14399
rect 31493 14365 31527 14399
rect 31585 14365 31619 14399
rect 31769 14365 31803 14399
rect 1685 14297 1719 14331
rect 5917 14297 5951 14331
rect 9597 14297 9631 14331
rect 19257 14297 19291 14331
rect 30573 14297 30607 14331
rect 30665 14297 30699 14331
rect 30849 14297 30883 14331
rect 13093 14229 13127 14263
rect 19634 14229 19668 14263
rect 31033 14229 31067 14263
rect 1961 14025 1995 14059
rect 6377 14025 6411 14059
rect 6653 14025 6687 14059
rect 7021 14025 7055 14059
rect 8677 14025 8711 14059
rect 17785 14025 17819 14059
rect 17877 14025 17911 14059
rect 19809 14025 19843 14059
rect 22845 14025 22879 14059
rect 23489 14025 23523 14059
rect 29101 14025 29135 14059
rect 31401 14025 31435 14059
rect 32873 14025 32907 14059
rect 7113 13957 7147 13991
rect 17233 13957 17267 13991
rect 25421 13957 25455 13991
rect 26433 13957 26467 13991
rect 1777 13889 1811 13923
rect 2145 13889 2179 13923
rect 6561 13889 6595 13923
rect 8401 13889 8435 13923
rect 8493 13889 8527 13923
rect 14657 13889 14691 13923
rect 15301 13889 15335 13923
rect 16221 13889 16255 13923
rect 16681 13889 16715 13923
rect 16773 13889 16807 13923
rect 19717 13889 19751 13923
rect 20269 13889 20303 13923
rect 20637 13889 20671 13923
rect 20913 13889 20947 13923
rect 21097 13889 21131 13923
rect 21189 13889 21223 13923
rect 21282 13879 21316 13913
rect 22109 13889 22143 13923
rect 22293 13889 22327 13923
rect 22661 13889 22695 13923
rect 24133 13889 24167 13923
rect 24409 13889 24443 13923
rect 24777 13889 24811 13923
rect 24869 13889 24903 13923
rect 25053 13889 25087 13923
rect 25145 13889 25179 13923
rect 25605 13889 25639 13923
rect 25697 13889 25731 13923
rect 25881 13889 25915 13923
rect 25973 13889 26007 13923
rect 26065 13889 26099 13923
rect 26249 13889 26283 13923
rect 26341 13889 26375 13923
rect 26525 13889 26559 13923
rect 26617 13889 26651 13923
rect 26801 13889 26835 13923
rect 27077 13889 27111 13923
rect 27261 13889 27295 13923
rect 28825 13889 28859 13923
rect 29101 13889 29135 13923
rect 29285 13889 29319 13923
rect 30205 13889 30239 13923
rect 30389 13889 30423 13923
rect 30757 13889 30791 13923
rect 30941 13889 30975 13923
rect 31953 13889 31987 13923
rect 32781 13889 32815 13923
rect 32965 13889 32999 13923
rect 33057 13889 33091 13923
rect 33241 13889 33275 13923
rect 1501 13821 1535 13855
rect 7205 13821 7239 13855
rect 15577 13821 15611 13855
rect 17969 13821 18003 13855
rect 21925 13821 21959 13855
rect 22477 13821 22511 13855
rect 23029 13821 23063 13855
rect 23121 13821 23155 13855
rect 23213 13821 23247 13855
rect 23305 13821 23339 13855
rect 23673 13821 23707 13855
rect 28917 13821 28951 13855
rect 30481 13821 30515 13855
rect 30573 13821 30607 13855
rect 31677 13821 31711 13855
rect 21557 13753 21591 13787
rect 24409 13753 24443 13787
rect 25329 13753 25363 13787
rect 15025 13685 15059 13719
rect 17417 13685 17451 13719
rect 26157 13685 26191 13719
rect 26801 13685 26835 13719
rect 27169 13685 27203 13719
rect 28549 13685 28583 13719
rect 31861 13685 31895 13719
rect 33241 13685 33275 13719
rect 4261 13481 4295 13515
rect 10517 13481 10551 13515
rect 15393 13481 15427 13515
rect 16681 13481 16715 13515
rect 17877 13481 17911 13515
rect 18429 13481 18463 13515
rect 18889 13481 18923 13515
rect 19717 13481 19751 13515
rect 20637 13481 20671 13515
rect 27445 13481 27479 13515
rect 28089 13481 28123 13515
rect 29101 13481 29135 13515
rect 29193 13481 29227 13515
rect 33149 13481 33183 13515
rect 33241 13481 33275 13515
rect 33701 13481 33735 13515
rect 9137 13413 9171 13447
rect 18613 13413 18647 13447
rect 20821 13413 20855 13447
rect 22661 13413 22695 13447
rect 22937 13413 22971 13447
rect 28273 13413 28307 13447
rect 4353 13345 4387 13379
rect 6377 13345 6411 13379
rect 7205 13345 7239 13379
rect 9781 13345 9815 13379
rect 10977 13345 11011 13379
rect 12909 13345 12943 13379
rect 13093 13345 13127 13379
rect 26249 13345 26283 13379
rect 26341 13345 26375 13379
rect 26709 13345 26743 13379
rect 29009 13345 29043 13379
rect 32965 13345 32999 13379
rect 34069 13345 34103 13379
rect 3893 13277 3927 13311
rect 8769 13277 8803 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 10609 13277 10643 13311
rect 10701 13277 10735 13311
rect 13185 13277 13219 13311
rect 13829 13277 13863 13311
rect 17785 13277 17819 13311
rect 19993 13277 20027 13311
rect 20085 13277 20119 13311
rect 20177 13277 20211 13311
rect 20361 13277 20395 13311
rect 21097 13277 21131 13311
rect 21373 13277 21407 13311
rect 21741 13277 21775 13311
rect 22385 13277 22419 13311
rect 22569 13277 22603 13311
rect 22937 13277 22971 13311
rect 23213 13277 23247 13311
rect 23489 13277 23523 13311
rect 24409 13277 24443 13311
rect 24685 13277 24719 13311
rect 25697 13277 25731 13311
rect 25881 13277 25915 13311
rect 25973 13277 26007 13311
rect 26157 13277 26191 13311
rect 26525 13277 26559 13311
rect 26801 13277 26835 13311
rect 26985 13277 27019 13311
rect 27077 13277 27111 13311
rect 27169 13277 27203 13311
rect 28365 13277 28399 13311
rect 28457 13277 28491 13311
rect 28549 13277 28583 13311
rect 28733 13277 28767 13311
rect 29285 13277 29319 13311
rect 29561 13277 29595 13311
rect 29745 13277 29779 13311
rect 32873 13277 32907 13311
rect 33425 13277 33459 13311
rect 33517 13277 33551 13311
rect 33885 13277 33919 13311
rect 18843 13243 18877 13277
rect 4077 13209 4111 13243
rect 4629 13209 4663 13243
rect 6929 13209 6963 13243
rect 9965 13209 9999 13243
rect 11253 13209 11287 13243
rect 15025 13209 15059 13243
rect 15209 13209 15243 13243
rect 16681 13209 16715 13243
rect 16865 13209 16899 13243
rect 18245 13209 18279 13243
rect 19073 13209 19107 13243
rect 20453 13209 20487 13243
rect 20653 13209 20687 13243
rect 21005 13209 21039 13243
rect 23305 13209 23339 13243
rect 23673 13209 23707 13243
rect 24777 13209 24811 13243
rect 32505 13209 32539 13243
rect 32597 13209 32631 13243
rect 6561 13141 6595 13175
rect 7021 13141 7055 13175
rect 8585 13141 8619 13175
rect 9505 13141 9539 13175
rect 9597 13141 9631 13175
rect 10885 13141 10919 13175
rect 12725 13141 12759 13175
rect 13553 13141 13587 13175
rect 13645 13141 13679 13175
rect 16497 13141 16531 13175
rect 18445 13141 18479 13175
rect 18705 13141 18739 13175
rect 21557 13141 21591 13175
rect 25789 13141 25823 13175
rect 29653 13141 29687 13175
rect 3157 12937 3191 12971
rect 4997 12937 5031 12971
rect 8125 12937 8159 12971
rect 14933 12937 14967 12971
rect 19743 12937 19777 12971
rect 20361 12937 20395 12971
rect 21649 12937 21683 12971
rect 24869 12937 24903 12971
rect 26249 12937 26283 12971
rect 31217 12937 31251 12971
rect 31861 12937 31895 12971
rect 32873 12937 32907 12971
rect 4077 12869 4111 12903
rect 4537 12869 4571 12903
rect 8585 12869 8619 12903
rect 13461 12869 13495 12903
rect 19533 12869 19567 12903
rect 31493 12869 31527 12903
rect 31709 12869 31743 12903
rect 32505 12869 32539 12903
rect 1409 12801 1443 12835
rect 3985 12801 4019 12835
rect 4445 12801 4479 12835
rect 4629 12801 4663 12835
rect 5181 12801 5215 12835
rect 6009 12801 6043 12835
rect 6377 12801 6411 12835
rect 8309 12801 8343 12835
rect 10333 12801 10367 12835
rect 10517 12801 10551 12835
rect 10609 12801 10643 12835
rect 13093 12801 13127 12835
rect 15485 12801 15519 12835
rect 16865 12801 16899 12835
rect 20177 12801 20211 12835
rect 20545 12801 20579 12835
rect 21097 12801 21131 12835
rect 21465 12801 21499 12835
rect 21833 12801 21867 12835
rect 24961 12801 24995 12835
rect 25053 12801 25087 12835
rect 26433 12801 26467 12835
rect 26525 12801 26559 12835
rect 26709 12801 26743 12835
rect 26801 12801 26835 12835
rect 29101 12801 29135 12835
rect 30665 12801 30699 12835
rect 31217 12801 31251 12835
rect 31401 12801 31435 12835
rect 32137 12801 32171 12835
rect 32321 12801 32355 12835
rect 33149 12801 33183 12835
rect 1685 12733 1719 12767
rect 4169 12733 4203 12767
rect 6653 12733 6687 12767
rect 12265 12733 12299 12767
rect 13185 12733 13219 12767
rect 15577 12733 15611 12767
rect 15669 12733 15703 12767
rect 17601 12733 17635 12767
rect 22201 12733 22235 12767
rect 22293 12733 22327 12767
rect 22385 12733 22419 12767
rect 24409 12733 24443 12767
rect 24501 12733 24535 12767
rect 24593 12733 24627 12767
rect 24685 12733 24719 12767
rect 25237 12733 25271 12767
rect 29377 12733 29411 12767
rect 30573 12733 30607 12767
rect 32873 12733 32907 12767
rect 33057 12733 33091 12767
rect 6193 12665 6227 12699
rect 10057 12665 10091 12699
rect 29193 12665 29227 12699
rect 31033 12665 31067 12699
rect 3617 12597 3651 12631
rect 10149 12597 10183 12631
rect 15117 12597 15151 12631
rect 19717 12597 19751 12631
rect 19901 12597 19935 12631
rect 20177 12597 20211 12631
rect 21465 12597 21499 12631
rect 25145 12597 25179 12631
rect 29285 12597 29319 12631
rect 31677 12597 31711 12631
rect 1961 12393 1995 12427
rect 3801 12393 3835 12427
rect 3985 12393 4019 12427
rect 4261 12393 4295 12427
rect 6469 12393 6503 12427
rect 8585 12393 8619 12427
rect 11529 12393 11563 12427
rect 14933 12393 14967 12427
rect 15374 12393 15408 12427
rect 16865 12393 16899 12427
rect 21741 12393 21775 12427
rect 25237 12393 25271 12427
rect 26893 12393 26927 12427
rect 29561 12393 29595 12427
rect 30205 12393 30239 12427
rect 23673 12325 23707 12359
rect 3065 12257 3099 12291
rect 3249 12257 3283 12291
rect 6929 12257 6963 12291
rect 7113 12257 7147 12291
rect 11989 12257 12023 12291
rect 12173 12257 12207 12291
rect 18153 12257 18187 12291
rect 18429 12257 18463 12291
rect 22937 12257 22971 12291
rect 23029 12257 23063 12291
rect 23121 12257 23155 12291
rect 23581 12257 23615 12291
rect 23765 12257 23799 12291
rect 25789 12257 25823 12291
rect 26249 12257 26283 12291
rect 30297 12257 30331 12291
rect 2145 12189 2179 12223
rect 2973 12189 3007 12223
rect 4261 12189 4295 12223
rect 4537 12189 4571 12223
rect 8217 12189 8251 12223
rect 8401 12189 8435 12223
rect 9965 12189 9999 12223
rect 10149 12189 10183 12223
rect 14749 12189 14783 12223
rect 15117 12189 15151 12223
rect 18613 12189 18647 12223
rect 18981 12189 19015 12223
rect 19349 12189 19383 12223
rect 23213 12189 23247 12223
rect 23489 12189 23523 12223
rect 25605 12189 25639 12223
rect 26433 12189 26467 12223
rect 29837 12189 29871 12223
rect 30021 12189 30055 12223
rect 30389 12189 30423 12223
rect 30573 12189 30607 12223
rect 33149 12189 33183 12223
rect 33517 12189 33551 12223
rect 4169 12121 4203 12155
rect 4445 12121 4479 12155
rect 6837 12121 6871 12155
rect 8677 12121 8711 12155
rect 11897 12121 11931 12155
rect 18061 12121 18095 12155
rect 18889 12121 18923 12155
rect 21557 12121 21591 12155
rect 21773 12121 21807 12155
rect 29929 12121 29963 12155
rect 2605 12053 2639 12087
rect 3959 12053 3993 12087
rect 8033 12053 8067 12087
rect 9781 12053 9815 12087
rect 17601 12053 17635 12087
rect 17969 12053 18003 12087
rect 19533 12053 19567 12087
rect 21925 12053 21959 12087
rect 23397 12053 23431 12087
rect 25697 12053 25731 12087
rect 26525 12053 26559 12087
rect 30481 12053 30515 12087
rect 33149 12053 33183 12087
rect 24402 11849 24436 11883
rect 29285 11849 29319 11883
rect 29745 11849 29779 11883
rect 32413 11849 32447 11883
rect 12541 11781 12575 11815
rect 27905 11781 27939 11815
rect 30205 11781 30239 11815
rect 1501 11713 1535 11747
rect 1685 11713 1719 11747
rect 10701 11713 10735 11747
rect 10793 11713 10827 11747
rect 11989 11713 12023 11747
rect 15945 11713 15979 11747
rect 18613 11713 18647 11747
rect 18797 11713 18831 11747
rect 23581 11713 23615 11747
rect 23765 11713 23799 11747
rect 24225 11713 24259 11747
rect 24317 11713 24351 11747
rect 24501 11713 24535 11747
rect 24593 11713 24627 11747
rect 24777 11713 24811 11747
rect 24869 11713 24903 11747
rect 25053 11713 25087 11747
rect 27169 11713 27203 11747
rect 27353 11713 27387 11747
rect 27442 11735 27476 11769
rect 27675 11747 27709 11781
rect 29469 11713 29503 11747
rect 29929 11713 29963 11747
rect 30573 11713 30607 11747
rect 32597 11713 32631 11747
rect 32689 11713 32723 11747
rect 10885 11645 10919 11679
rect 12265 11645 12299 11679
rect 14289 11645 14323 11679
rect 16037 11645 16071 11679
rect 16129 11645 16163 11679
rect 24961 11645 24995 11679
rect 29561 11645 29595 11679
rect 29837 11645 29871 11679
rect 30665 11645 30699 11679
rect 12173 11577 12207 11611
rect 18705 11577 18739 11611
rect 24593 11577 24627 11611
rect 27537 11577 27571 11611
rect 10333 11509 10367 11543
rect 15577 11509 15611 11543
rect 23581 11509 23615 11543
rect 26985 11509 27019 11543
rect 27721 11509 27755 11543
rect 30849 11509 30883 11543
rect 3157 11305 3191 11339
rect 5733 11305 5767 11339
rect 8493 11305 8527 11339
rect 12449 11305 12483 11339
rect 17601 11305 17635 11339
rect 28917 11305 28951 11339
rect 29285 11305 29319 11339
rect 31401 11305 31435 11339
rect 32137 11305 32171 11339
rect 8033 11237 8067 11271
rect 9321 11237 9355 11271
rect 9965 11237 9999 11271
rect 14105 11237 14139 11271
rect 15761 11237 15795 11271
rect 21925 11237 21959 11271
rect 30573 11237 30607 11271
rect 1409 11169 1443 11203
rect 4353 11169 4387 11203
rect 8309 11169 8343 11203
rect 9229 11169 9263 11203
rect 10057 11169 10091 11203
rect 10333 11169 10367 11203
rect 11805 11169 11839 11203
rect 12909 11169 12943 11203
rect 13093 11169 13127 11203
rect 14749 11169 14783 11203
rect 16129 11169 16163 11203
rect 23765 11169 23799 11203
rect 26157 11169 26191 11203
rect 27169 11169 27203 11203
rect 30113 11169 30147 11203
rect 5917 11101 5951 11135
rect 6101 11101 6135 11135
rect 7389 11101 7423 11135
rect 7481 11101 7515 11135
rect 7665 11101 7699 11135
rect 7757 11101 7791 11135
rect 8585 11101 8619 11135
rect 9137 11101 9171 11135
rect 9413 11101 9447 11135
rect 9781 11101 9815 11135
rect 13737 11101 13771 11135
rect 14473 11101 14507 11135
rect 15577 11101 15611 11135
rect 15853 11101 15887 11135
rect 18613 11101 18647 11135
rect 18797 11101 18831 11135
rect 19257 11101 19291 11135
rect 19901 11101 19935 11135
rect 19993 11101 20027 11135
rect 20085 11101 20119 11135
rect 21373 11101 21407 11135
rect 21649 11101 21683 11135
rect 21741 11101 21775 11135
rect 22017 11101 22051 11135
rect 22201 11101 22235 11135
rect 22477 11101 22511 11135
rect 23581 11101 23615 11135
rect 25421 11101 25455 11135
rect 25605 11101 25639 11135
rect 26433 11101 26467 11135
rect 26893 11101 26927 11135
rect 27077 11101 27111 11135
rect 27261 11101 27295 11135
rect 27445 11101 27479 11135
rect 27721 11101 27755 11135
rect 27905 11101 27939 11135
rect 28181 11101 28215 11135
rect 28273 11101 28307 11135
rect 28457 11101 28491 11135
rect 29101 11101 29135 11135
rect 29377 11101 29411 11135
rect 30205 11101 30239 11135
rect 30297 11101 30331 11135
rect 30389 11101 30423 11135
rect 31585 11101 31619 11135
rect 31861 11101 31895 11135
rect 32045 11101 32079 11135
rect 32321 11101 32355 11135
rect 32597 11101 32631 11135
rect 32781 11101 32815 11135
rect 32873 11101 32907 11135
rect 33057 11101 33091 11135
rect 37565 11101 37599 11135
rect 1685 11033 1719 11067
rect 4169 11033 4203 11067
rect 7941 11033 7975 11067
rect 8953 11033 8987 11067
rect 12817 11033 12851 11067
rect 18429 11033 18463 11067
rect 19533 11033 19567 11067
rect 20269 11033 20303 11067
rect 21557 11033 21591 11067
rect 22385 11033 22419 11067
rect 25513 11033 25547 11067
rect 28089 11033 28123 11067
rect 37933 11033 37967 11067
rect 3801 10965 3835 10999
rect 4261 10965 4295 10999
rect 13921 10965 13955 10999
rect 14565 10965 14599 10999
rect 23397 10965 23431 10999
rect 26341 10965 26375 10999
rect 26801 10965 26835 10999
rect 27629 10965 27663 10999
rect 28457 10965 28491 10999
rect 32965 10965 32999 10999
rect 1777 10761 1811 10795
rect 2789 10761 2823 10795
rect 5825 10761 5859 10795
rect 8677 10761 8711 10795
rect 9045 10761 9079 10795
rect 19165 10761 19199 10795
rect 24133 10761 24167 10795
rect 24225 10761 24259 10795
rect 32229 10761 32263 10795
rect 33701 10761 33735 10795
rect 35081 10761 35115 10795
rect 7389 10693 7423 10727
rect 7573 10693 7607 10727
rect 14197 10693 14231 10727
rect 15945 10693 15979 10727
rect 20821 10693 20855 10727
rect 21021 10693 21055 10727
rect 23121 10693 23155 10727
rect 23259 10693 23293 10727
rect 28549 10693 28583 10727
rect 1961 10625 1995 10659
rect 2697 10625 2731 10659
rect 3341 10625 3375 10659
rect 6009 10625 6043 10659
rect 6193 10625 6227 10659
rect 6745 10625 6779 10659
rect 7205 10625 7239 10659
rect 8585 10625 8619 10659
rect 8861 10625 8895 10659
rect 9597 10625 9631 10659
rect 10977 10625 11011 10659
rect 13921 10625 13955 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 17141 10625 17175 10659
rect 17233 10625 17267 10659
rect 18153 10625 18187 10659
rect 18337 10625 18371 10659
rect 18981 10625 19015 10659
rect 20269 10625 20303 10659
rect 21465 10625 21499 10659
rect 22109 10625 22143 10659
rect 22201 10625 22235 10659
rect 22385 10625 22419 10659
rect 22477 10625 22511 10659
rect 22938 10647 22972 10681
rect 23029 10625 23063 10659
rect 26985 10625 27019 10659
rect 27169 10625 27203 10659
rect 27261 10625 27295 10659
rect 27353 10625 27387 10659
rect 28273 10625 28307 10659
rect 28365 10625 28399 10659
rect 28733 10625 28767 10659
rect 28917 10625 28951 10659
rect 30297 10625 30331 10659
rect 30481 10625 30515 10659
rect 32137 10625 32171 10659
rect 32321 10625 32355 10659
rect 32597 10625 32631 10659
rect 33517 10625 33551 10659
rect 33793 10625 33827 10659
rect 34069 10625 34103 10659
rect 34713 10625 34747 10659
rect 2973 10557 3007 10591
rect 3433 10557 3467 10591
rect 3709 10557 3743 10591
rect 4077 10557 4111 10591
rect 4353 10557 4387 10591
rect 6101 10557 6135 10591
rect 6837 10557 6871 10591
rect 6929 10557 6963 10591
rect 9137 10557 9171 10591
rect 11069 10557 11103 10591
rect 11253 10557 11287 10591
rect 21281 10557 21315 10591
rect 21649 10557 21683 10591
rect 21925 10557 21959 10591
rect 23397 10557 23431 10591
rect 23949 10557 23983 10591
rect 30389 10557 30423 10591
rect 32505 10557 32539 10591
rect 33977 10557 34011 10591
rect 34621 10557 34655 10591
rect 2329 10489 2363 10523
rect 17509 10489 17543 10523
rect 24593 10489 24627 10523
rect 28733 10489 28767 10523
rect 34437 10489 34471 10523
rect 6377 10421 6411 10455
rect 9321 10421 9355 10455
rect 10609 10421 10643 10455
rect 18061 10421 18095 10455
rect 20177 10421 20211 10455
rect 21005 10421 21039 10455
rect 21189 10421 21223 10455
rect 22753 10421 22787 10455
rect 27629 10421 27663 10455
rect 32873 10421 32907 10455
rect 33517 10421 33551 10455
rect 4629 10217 4663 10251
rect 6193 10217 6227 10251
rect 7573 10217 7607 10251
rect 20453 10217 20487 10251
rect 20913 10217 20947 10251
rect 22385 10217 22419 10251
rect 22661 10217 22695 10251
rect 32689 10217 32723 10251
rect 33517 10217 33551 10251
rect 8493 10149 8527 10183
rect 20821 10149 20855 10183
rect 21189 10149 21223 10183
rect 21649 10149 21683 10183
rect 29009 10149 29043 10183
rect 5641 10081 5675 10115
rect 5825 10081 5859 10115
rect 7757 10081 7791 10115
rect 8334 10081 8368 10115
rect 9045 10081 9079 10115
rect 9321 10081 9355 10115
rect 11713 10081 11747 10115
rect 17601 10081 17635 10115
rect 21281 10081 21315 10115
rect 21373 10081 21407 10115
rect 22385 10081 22419 10115
rect 30389 10081 30423 10115
rect 30481 10081 30515 10115
rect 2973 10013 3007 10047
rect 4813 10013 4847 10047
rect 5549 10013 5583 10047
rect 6009 10013 6043 10047
rect 6193 10013 6227 10047
rect 7481 10013 7515 10047
rect 7849 10013 7883 10047
rect 9137 10013 9171 10047
rect 9229 10013 9263 10047
rect 11437 10013 11471 10047
rect 13737 10013 13771 10047
rect 17785 10013 17819 10047
rect 18061 10013 18095 10047
rect 18245 10013 18279 10047
rect 18337 10013 18371 10047
rect 18429 10013 18463 10047
rect 20269 10013 20303 10047
rect 20453 10013 20487 10047
rect 20545 10013 20579 10047
rect 21097 10013 21131 10047
rect 21557 10013 21591 10047
rect 21649 10013 21683 10047
rect 21833 10013 21867 10047
rect 21925 10013 21959 10047
rect 22293 10013 22327 10047
rect 28273 10013 28307 10047
rect 28641 10013 28675 10047
rect 28733 10013 28767 10047
rect 28917 10013 28951 10047
rect 30113 10013 30147 10047
rect 30297 10013 30331 10047
rect 30665 10013 30699 10047
rect 32597 10013 32631 10047
rect 33793 10013 33827 10047
rect 33885 10013 33919 10047
rect 33977 10013 34011 10047
rect 34161 10013 34195 10047
rect 2789 9945 2823 9979
rect 11989 9945 12023 9979
rect 17969 9945 18003 9979
rect 19349 9945 19383 9979
rect 19717 9945 19751 9979
rect 20637 9945 20671 9979
rect 20821 9945 20855 9979
rect 28457 9945 28491 9979
rect 3157 9877 3191 9911
rect 5181 9877 5215 9911
rect 7757 9877 7791 9911
rect 8125 9877 8159 9911
rect 8217 9877 8251 9911
rect 9505 9877 9539 9911
rect 11621 9877 11655 9911
rect 18705 9877 18739 9911
rect 30849 9877 30883 9911
rect 11805 9673 11839 9707
rect 13093 9673 13127 9707
rect 13461 9673 13495 9707
rect 15945 9673 15979 9707
rect 22477 9673 22511 9707
rect 33241 9673 33275 9707
rect 6377 9605 6411 9639
rect 8309 9605 8343 9639
rect 8585 9605 8619 9639
rect 10793 9605 10827 9639
rect 15485 9605 15519 9639
rect 23121 9605 23155 9639
rect 24593 9605 24627 9639
rect 24685 9605 24719 9639
rect 26341 9605 26375 9639
rect 30021 9605 30055 9639
rect 33057 9605 33091 9639
rect 3249 9537 3283 9571
rect 3341 9537 3375 9571
rect 3433 9537 3467 9571
rect 3617 9537 3651 9571
rect 6653 9537 6687 9571
rect 6745 9537 6779 9571
rect 6837 9537 6871 9571
rect 7021 9537 7055 9571
rect 7757 9537 7791 9571
rect 8033 9537 8067 9571
rect 8493 9537 8527 9571
rect 8677 9537 8711 9571
rect 10241 9537 10275 9571
rect 10701 9537 10735 9571
rect 12173 9537 12207 9571
rect 12265 9537 12299 9571
rect 15577 9537 15611 9571
rect 16221 9537 16255 9571
rect 16773 9537 16807 9571
rect 18429 9537 18463 9571
rect 18797 9537 18831 9571
rect 19809 9537 19843 9571
rect 19901 9537 19935 9571
rect 20085 9537 20119 9571
rect 22661 9537 22695 9571
rect 22753 9537 22787 9571
rect 23029 9537 23063 9571
rect 24133 9537 24167 9571
rect 24317 9537 24351 9571
rect 24409 9537 24443 9571
rect 24777 9537 24811 9571
rect 25973 9537 26007 9571
rect 26157 9537 26191 9571
rect 26433 9537 26467 9571
rect 26617 9537 26651 9571
rect 26985 9537 27019 9571
rect 27169 9537 27203 9571
rect 27445 9537 27479 9571
rect 28825 9537 28859 9571
rect 29009 9537 29043 9571
rect 29653 9537 29687 9571
rect 29745 9537 29779 9571
rect 29837 9537 29871 9571
rect 29929 9537 29963 9571
rect 30113 9537 30147 9571
rect 30757 9537 30791 9571
rect 31033 9537 31067 9571
rect 31309 9537 31343 9571
rect 31585 9537 31619 9571
rect 32505 9537 32539 9571
rect 32873 9537 32907 9571
rect 10885 9469 10919 9503
rect 12449 9469 12483 9503
rect 13553 9469 13587 9503
rect 13645 9469 13679 9503
rect 15301 9469 15335 9503
rect 17233 9469 17267 9503
rect 18245 9469 18279 9503
rect 18705 9469 18739 9503
rect 19441 9469 19475 9503
rect 19993 9469 20027 9503
rect 32413 9469 32447 9503
rect 7481 9401 7515 9435
rect 8033 9401 8067 9435
rect 10333 9401 10367 9435
rect 24317 9401 24351 9435
rect 24961 9401 24995 9435
rect 31217 9401 31251 9435
rect 32137 9401 32171 9435
rect 2973 9333 3007 9367
rect 10057 9333 10091 9367
rect 16037 9333 16071 9367
rect 19625 9333 19659 9367
rect 26525 9333 26559 9367
rect 27629 9333 27663 9367
rect 29193 9333 29227 9367
rect 6193 9129 6227 9163
rect 11529 9129 11563 9163
rect 17509 9129 17543 9163
rect 20913 9129 20947 9163
rect 23949 9129 23983 9163
rect 29745 9129 29779 9163
rect 31769 9129 31803 9163
rect 32873 9129 32907 9163
rect 33241 9129 33275 9163
rect 22845 9061 22879 9095
rect 29929 9061 29963 9095
rect 32413 9061 32447 9095
rect 4629 8993 4663 9027
rect 8677 8993 8711 9027
rect 9781 8993 9815 9027
rect 10057 8993 10091 9027
rect 13645 8993 13679 9027
rect 15577 8993 15611 9027
rect 18337 8993 18371 9027
rect 20269 8993 20303 9027
rect 20729 8993 20763 9027
rect 22201 8993 22235 9027
rect 22661 8993 22695 9027
rect 25329 8993 25363 9027
rect 25789 8993 25823 9027
rect 27077 8993 27111 9027
rect 29285 8993 29319 9027
rect 31493 8993 31527 9027
rect 33517 8993 33551 9027
rect 1777 8925 1811 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 4353 8925 4387 8959
rect 4537 8925 4571 8959
rect 4997 8925 5031 8959
rect 5825 8925 5859 8959
rect 12725 8925 12759 8959
rect 12909 8925 12943 8959
rect 13369 8925 13403 8959
rect 14093 8925 14127 8959
rect 14289 8925 14323 8959
rect 14384 8925 14418 8959
rect 14519 8925 14553 8959
rect 15301 8925 15335 8959
rect 15761 8925 15795 8959
rect 17969 8925 18003 8959
rect 18705 8925 18739 8959
rect 19717 8925 19751 8959
rect 19901 8925 19935 8959
rect 19993 8925 20027 8959
rect 20637 8925 20671 8959
rect 22569 8925 22603 8959
rect 22937 8925 22971 8959
rect 23030 8925 23064 8959
rect 23213 8925 23247 8959
rect 23402 8925 23436 8959
rect 23857 8925 23891 8959
rect 24409 8925 24443 8959
rect 24502 8925 24536 8959
rect 24685 8925 24719 8959
rect 24777 8925 24811 8959
rect 24915 8925 24949 8959
rect 25237 8925 25271 8959
rect 25513 8925 25547 8959
rect 25605 8925 25639 8959
rect 25881 8925 25915 8959
rect 26065 8925 26099 8959
rect 26157 8925 26191 8959
rect 26249 8925 26283 8959
rect 26801 8925 26835 8959
rect 26985 8925 27019 8959
rect 27169 8925 27203 8959
rect 27353 8925 27387 8959
rect 27629 8925 27663 8959
rect 27997 8925 28031 8959
rect 28181 8925 28215 8959
rect 28365 8925 28399 8959
rect 28457 8925 28491 8959
rect 28549 8925 28583 8959
rect 28917 8925 28951 8959
rect 29101 8925 29135 8959
rect 29199 8925 29233 8959
rect 29377 8925 29411 8959
rect 29561 8925 29595 8959
rect 29653 8925 29687 8959
rect 30021 8925 30055 8959
rect 30205 8925 30239 8959
rect 31585 8925 31619 8959
rect 31861 8925 31895 8959
rect 32137 8925 32171 8959
rect 32597 8925 32631 8959
rect 32689 8925 32723 8959
rect 32965 8925 32999 8959
rect 33057 8925 33091 8959
rect 33241 8925 33275 8959
rect 37933 8925 37967 8959
rect 1409 8857 1443 8891
rect 4813 8857 4847 8891
rect 6009 8857 6043 8891
rect 12817 8857 12851 8891
rect 15393 8857 15427 8891
rect 16037 8857 16071 8891
rect 19533 8857 19567 8891
rect 22293 8857 22327 8891
rect 23305 8857 23339 8891
rect 27813 8857 27847 8891
rect 30389 8857 30423 8891
rect 37657 8857 37691 8891
rect 3893 8789 3927 8823
rect 8033 8789 8067 8823
rect 8401 8789 8435 8823
rect 8493 8789 8527 8823
rect 13001 8789 13035 8823
rect 13461 8789 13495 8823
rect 14749 8789 14783 8823
rect 14933 8789 14967 8823
rect 23581 8789 23615 8823
rect 25053 8789 25087 8823
rect 26525 8789 26559 8823
rect 27537 8789 27571 8823
rect 28825 8789 28859 8823
rect 29009 8789 29043 8823
rect 31125 8789 31159 8823
rect 31953 8789 31987 8823
rect 4261 8585 4295 8619
rect 5089 8585 5123 8619
rect 6377 8585 6411 8619
rect 9689 8585 9723 8619
rect 10057 8585 10091 8619
rect 10609 8585 10643 8619
rect 15209 8585 15243 8619
rect 18889 8585 18923 8619
rect 24961 8585 24995 8619
rect 29285 8585 29319 8619
rect 31309 8585 31343 8619
rect 6529 8517 6563 8551
rect 6745 8517 6779 8551
rect 7849 8517 7883 8551
rect 12449 8517 12483 8551
rect 12633 8517 12667 8551
rect 19533 8517 19567 8551
rect 22109 8517 22143 8551
rect 3433 8449 3467 8483
rect 4169 8449 4203 8483
rect 5457 8449 5491 8483
rect 5917 8449 5951 8483
rect 6101 8449 6135 8483
rect 6193 8449 6227 8483
rect 9597 8449 9631 8483
rect 10149 8449 10183 8483
rect 10517 8449 10551 8483
rect 11529 8449 11563 8483
rect 11989 8449 12023 8483
rect 12357 8449 12391 8483
rect 12541 8449 12575 8483
rect 13001 8449 13035 8483
rect 13185 8449 13219 8483
rect 13461 8449 13495 8483
rect 17417 8449 17451 8483
rect 17509 8449 17543 8483
rect 18797 8449 18831 8483
rect 18981 8449 19015 8483
rect 19717 8449 19751 8483
rect 19809 8449 19843 8483
rect 21925 8449 21959 8483
rect 23213 8449 23247 8483
rect 23489 8449 23523 8483
rect 23673 8449 23707 8483
rect 24869 8449 24903 8483
rect 26985 8449 27019 8483
rect 27169 8449 27203 8483
rect 27261 8449 27295 8483
rect 27353 8449 27387 8483
rect 27537 8449 27571 8483
rect 28917 8449 28951 8483
rect 29101 8449 29135 8483
rect 31585 8449 31619 8483
rect 31861 8449 31895 8483
rect 33149 8449 33183 8483
rect 4445 8381 4479 8415
rect 5549 8381 5583 8415
rect 5641 8381 5675 8415
rect 10333 8381 10367 8415
rect 11897 8381 11931 8415
rect 13737 8381 13771 8415
rect 24777 8381 24811 8415
rect 31401 8381 31435 8415
rect 33241 8381 33275 8415
rect 3801 8313 3835 8347
rect 13369 8313 13403 8347
rect 17233 8313 17267 8347
rect 27721 8313 27755 8347
rect 32781 8313 32815 8347
rect 3249 8245 3283 8279
rect 5917 8245 5951 8279
rect 6561 8245 6595 8279
rect 19533 8245 19567 8279
rect 22293 8245 22327 8279
rect 23029 8245 23063 8279
rect 25329 8245 25363 8279
rect 29009 8245 29043 8279
rect 5641 8041 5675 8075
rect 8677 8041 8711 8075
rect 11897 8041 11931 8075
rect 12817 8041 12851 8075
rect 13553 8041 13587 8075
rect 13737 8041 13771 8075
rect 20177 8041 20211 8075
rect 31861 8041 31895 8075
rect 17509 7973 17543 8007
rect 21649 7973 21683 8007
rect 23305 7973 23339 8007
rect 30757 7973 30791 8007
rect 6653 7905 6687 7939
rect 6929 7905 6963 7939
rect 12633 7905 12667 7939
rect 15945 7905 15979 7939
rect 22385 7905 22419 7939
rect 30297 7905 30331 7939
rect 5641 7837 5675 7871
rect 5825 7837 5859 7871
rect 6469 7837 6503 7871
rect 9697 7837 9731 7871
rect 9873 7837 9907 7871
rect 10425 7837 10459 7871
rect 13369 7837 13403 7871
rect 13737 7837 13771 7871
rect 13921 7837 13955 7871
rect 15761 7837 15795 7871
rect 15853 7837 15887 7871
rect 17233 7837 17267 7871
rect 17601 7837 17635 7871
rect 17785 7837 17819 7871
rect 19717 7837 19751 7871
rect 19901 7837 19935 7871
rect 20085 7837 20119 7871
rect 20269 7837 20303 7871
rect 21557 7837 21591 7871
rect 21741 7837 21775 7871
rect 21833 7837 21867 7871
rect 21925 7837 21959 7871
rect 22109 7837 22143 7871
rect 22201 7837 22235 7871
rect 22661 7837 22695 7871
rect 30021 7837 30055 7871
rect 30205 7837 30239 7871
rect 30389 7837 30423 7871
rect 30573 7837 30607 7871
rect 30941 7837 30975 7871
rect 31401 7837 31435 7871
rect 31493 7837 31527 7871
rect 7205 7769 7239 7803
rect 12357 7769 12391 7803
rect 17509 7769 17543 7803
rect 17693 7769 17727 7803
rect 19809 7769 19843 7803
rect 22753 7769 22787 7803
rect 23121 7769 23155 7803
rect 31309 7769 31343 7803
rect 31677 7769 31711 7803
rect 6101 7701 6135 7735
rect 6561 7701 6595 7735
rect 9689 7701 9723 7735
rect 15393 7701 15427 7735
rect 17325 7701 17359 7735
rect 22293 7701 22327 7735
rect 31217 7701 31251 7735
rect 5641 7497 5675 7531
rect 7665 7497 7699 7531
rect 19625 7497 19659 7531
rect 22385 7497 22419 7531
rect 23213 7497 23247 7531
rect 26617 7497 26651 7531
rect 30113 7497 30147 7531
rect 2881 7429 2915 7463
rect 11805 7429 11839 7463
rect 19349 7429 19383 7463
rect 20177 7429 20211 7463
rect 22937 7429 22971 7463
rect 23949 7429 23983 7463
rect 25605 7429 25639 7463
rect 1501 7361 1535 7395
rect 2605 7361 2639 7395
rect 5549 7361 5583 7395
rect 6745 7361 6779 7395
rect 7849 7361 7883 7395
rect 14565 7361 14599 7395
rect 14841 7361 14875 7395
rect 15485 7361 15519 7395
rect 17785 7361 17819 7395
rect 17969 7361 18003 7395
rect 19165 7361 19199 7395
rect 19533 7361 19567 7395
rect 19809 7361 19843 7395
rect 20361 7361 20395 7395
rect 20821 7361 20855 7395
rect 21833 7361 21867 7395
rect 22109 7361 22143 7395
rect 22201 7361 22235 7395
rect 22569 7361 22603 7395
rect 22717 7361 22751 7395
rect 22845 7361 22879 7395
rect 23075 7361 23109 7395
rect 23857 7361 23891 7395
rect 24041 7361 24075 7395
rect 24133 7361 24167 7395
rect 24317 7361 24351 7395
rect 24501 7361 24535 7395
rect 24685 7361 24719 7395
rect 25145 7361 25179 7395
rect 26433 7361 26467 7395
rect 26617 7361 26651 7395
rect 27629 7361 27663 7395
rect 27813 7361 27847 7395
rect 27905 7361 27939 7395
rect 27997 7361 28031 7395
rect 28457 7361 28491 7395
rect 29009 7361 29043 7395
rect 29101 7361 29135 7395
rect 29377 7361 29411 7395
rect 29653 7361 29687 7395
rect 30113 7361 30147 7395
rect 30297 7361 30331 7395
rect 30757 7361 30791 7395
rect 31401 7361 31435 7395
rect 31769 7361 31803 7395
rect 31861 7361 31895 7395
rect 1685 7293 1719 7327
rect 4353 7293 4387 7327
rect 5825 7293 5859 7327
rect 6377 7293 6411 7327
rect 6837 7293 6871 7327
rect 9413 7293 9447 7327
rect 9689 7293 9723 7327
rect 11529 7293 11563 7327
rect 14473 7293 14507 7327
rect 14657 7293 14691 7327
rect 15025 7293 15059 7327
rect 18981 7293 19015 7327
rect 20913 7293 20947 7327
rect 24409 7293 24443 7327
rect 25329 7293 25363 7327
rect 27721 7293 27755 7327
rect 28273 7293 28307 7327
rect 31309 7293 31343 7327
rect 14197 7225 14231 7259
rect 19993 7225 20027 7259
rect 21189 7225 21223 7259
rect 5181 7157 5215 7191
rect 11161 7157 11195 7191
rect 13277 7157 13311 7191
rect 14565 7157 14599 7191
rect 15669 7157 15703 7191
rect 17877 7157 17911 7191
rect 21925 7157 21959 7191
rect 24869 7157 24903 7191
rect 24961 7157 24995 7191
rect 25145 7157 25179 7191
rect 6009 6953 6043 6987
rect 12357 6953 12391 6987
rect 12817 6953 12851 6987
rect 15742 6953 15776 6987
rect 17233 6953 17267 6987
rect 18061 6953 18095 6987
rect 25421 6953 25455 6987
rect 31493 6953 31527 6987
rect 17693 6885 17727 6919
rect 27077 6885 27111 6919
rect 30665 6885 30699 6919
rect 4261 6817 4295 6851
rect 12633 6817 12667 6851
rect 15485 6817 15519 6851
rect 17877 6817 17911 6851
rect 19993 6817 20027 6851
rect 20453 6817 20487 6851
rect 24869 6817 24903 6851
rect 27261 6817 27295 6851
rect 28549 6817 28583 6851
rect 32505 6817 32539 6851
rect 32597 6817 32631 6851
rect 32965 6817 32999 6851
rect 33149 6817 33183 6851
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 12909 6749 12943 6783
rect 15209 6749 15243 6783
rect 17601 6749 17635 6783
rect 17969 6749 18003 6783
rect 18153 6749 18187 6783
rect 18337 6749 18371 6783
rect 18429 6749 18463 6783
rect 18521 6749 18555 6783
rect 20085 6749 20119 6783
rect 21189 6749 21223 6783
rect 21281 6749 21315 6783
rect 21465 6749 21499 6783
rect 24961 6749 24995 6783
rect 25605 6749 25639 6783
rect 25697 6749 25731 6783
rect 25973 6749 26007 6783
rect 26157 6749 26191 6783
rect 26249 6749 26283 6783
rect 26341 6749 26375 6783
rect 26985 6749 27019 6783
rect 27537 6749 27571 6783
rect 27630 6749 27664 6783
rect 27905 6749 27939 6783
rect 28002 6749 28036 6783
rect 28273 6749 28307 6783
rect 28365 6749 28399 6783
rect 28733 6749 28767 6783
rect 29929 6749 29963 6783
rect 30113 6749 30147 6783
rect 30389 6749 30423 6783
rect 30757 6749 30791 6783
rect 30849 6749 30883 6783
rect 31769 6749 31803 6783
rect 31861 6749 31895 6783
rect 31953 6749 31987 6783
rect 32137 6749 32171 6783
rect 32689 6749 32723 6783
rect 32781 6749 32815 6783
rect 33241 6749 33275 6783
rect 4537 6681 4571 6715
rect 18797 6681 18831 6715
rect 25421 6681 25455 6715
rect 27261 6681 27295 6715
rect 27813 6681 27847 6715
rect 9045 6613 9079 6647
rect 14565 6613 14599 6647
rect 21649 6613 21683 6647
rect 25329 6613 25363 6647
rect 26617 6613 26651 6647
rect 28181 6613 28215 6647
rect 33609 6613 33643 6647
rect 4721 6409 4755 6443
rect 7849 6409 7883 6443
rect 14289 6409 14323 6443
rect 15301 6409 15335 6443
rect 18705 6409 18739 6443
rect 19901 6409 19935 6443
rect 23765 6409 23799 6443
rect 24231 6409 24265 6443
rect 25513 6409 25547 6443
rect 27997 6409 28031 6443
rect 28181 6409 28215 6443
rect 7757 6341 7791 6375
rect 9965 6341 9999 6375
rect 19073 6341 19107 6375
rect 22385 6341 22419 6375
rect 23397 6341 23431 6375
rect 23489 6341 23523 6375
rect 24133 6341 24167 6375
rect 32781 6341 32815 6375
rect 4905 6273 4939 6307
rect 8401 6273 8435 6307
rect 9505 6273 9539 6307
rect 9689 6273 9723 6307
rect 10057 6273 10091 6307
rect 12265 6273 12299 6307
rect 12449 6273 12483 6307
rect 12541 6273 12575 6307
rect 12817 6273 12851 6307
rect 13645 6273 13679 6307
rect 14565 6273 14599 6307
rect 15025 6273 15059 6307
rect 15393 6273 15427 6307
rect 15577 6273 15611 6307
rect 18061 6273 18095 6307
rect 18245 6273 18279 6307
rect 18337 6273 18371 6307
rect 18521 6273 18555 6307
rect 18889 6273 18923 6307
rect 19717 6273 19751 6307
rect 19901 6273 19935 6307
rect 22753 6273 22787 6307
rect 23213 6273 23247 6307
rect 23581 6273 23615 6307
rect 24317 6273 24351 6307
rect 24409 6273 24443 6307
rect 25421 6273 25455 6307
rect 25605 6273 25639 6307
rect 27813 6273 27847 6307
rect 28089 6273 28123 6307
rect 28273 6273 28307 6307
rect 32505 6273 32539 6307
rect 32597 6273 32631 6307
rect 7941 6205 7975 6239
rect 8585 6205 8619 6239
rect 8677 6205 8711 6239
rect 8769 6205 8803 6239
rect 9321 6205 9355 6239
rect 12081 6205 12115 6239
rect 14841 6205 14875 6239
rect 22845 6205 22879 6239
rect 27537 6205 27571 6239
rect 9689 6137 9723 6171
rect 18153 6137 18187 6171
rect 32781 6137 32815 6171
rect 7389 6069 7423 6103
rect 8217 6069 8251 6103
rect 15669 6069 15703 6103
rect 18521 6069 18555 6103
rect 19257 6069 19291 6103
rect 23029 6069 23063 6103
rect 27629 6069 27663 6103
rect 12817 5865 12851 5899
rect 15715 5865 15749 5899
rect 22661 5865 22695 5899
rect 30481 5865 30515 5899
rect 32045 5865 32079 5899
rect 32229 5865 32263 5899
rect 9137 5797 9171 5831
rect 22201 5797 22235 5831
rect 29837 5797 29871 5831
rect 5089 5729 5123 5763
rect 6929 5729 6963 5763
rect 7205 5729 7239 5763
rect 8677 5729 8711 5763
rect 9321 5729 9355 5763
rect 14933 5729 14967 5763
rect 17509 5729 17543 5763
rect 19257 5729 19291 5763
rect 19717 5729 19751 5763
rect 29561 5729 29595 5763
rect 9045 5661 9079 5695
rect 9413 5661 9447 5695
rect 9506 5661 9540 5695
rect 9781 5661 9815 5695
rect 9919 5661 9953 5695
rect 10149 5661 10183 5695
rect 10297 5661 10331 5695
rect 10655 5661 10689 5695
rect 12541 5661 12575 5695
rect 12725 5661 12759 5695
rect 12909 5661 12943 5695
rect 13645 5661 13679 5695
rect 13921 5661 13955 5695
rect 14749 5661 14783 5695
rect 15393 5661 15427 5695
rect 17141 5661 17175 5695
rect 19625 5661 19659 5695
rect 20085 5661 20119 5695
rect 20453 5661 20487 5695
rect 20637 5661 20671 5695
rect 22201 5661 22235 5695
rect 22385 5661 22419 5695
rect 22937 5661 22971 5695
rect 23121 5661 23155 5695
rect 23581 5661 23615 5695
rect 23673 5661 23707 5695
rect 24593 5661 24627 5695
rect 24869 5661 24903 5695
rect 25053 5661 25087 5695
rect 31861 5661 31895 5695
rect 32137 5661 32171 5695
rect 32321 5661 32355 5695
rect 5365 5593 5399 5627
rect 9689 5593 9723 5627
rect 10425 5593 10459 5627
rect 10517 5593 10551 5627
rect 11989 5593 12023 5627
rect 15485 5593 15519 5627
rect 19349 5593 19383 5627
rect 30113 5593 30147 5627
rect 30297 5593 30331 5627
rect 31677 5593 31711 5627
rect 6837 5525 6871 5559
rect 9045 5525 9079 5559
rect 10057 5525 10091 5559
rect 10793 5525 10827 5559
rect 13461 5525 13495 5559
rect 13829 5525 13863 5559
rect 14381 5525 14415 5559
rect 14841 5525 14875 5559
rect 19901 5525 19935 5559
rect 20453 5525 20487 5559
rect 24409 5525 24443 5559
rect 30021 5525 30055 5559
rect 6469 5321 6503 5355
rect 8861 5321 8895 5355
rect 15209 5321 15243 5355
rect 17325 5321 17359 5355
rect 19717 5321 19751 5355
rect 21281 5321 21315 5355
rect 23121 5321 23155 5355
rect 23673 5321 23707 5355
rect 27537 5321 27571 5355
rect 29469 5321 29503 5355
rect 30205 5321 30239 5355
rect 31493 5321 31527 5355
rect 9505 5253 9539 5287
rect 9689 5253 9723 5287
rect 11805 5253 11839 5287
rect 13737 5253 13771 5287
rect 19349 5253 19383 5287
rect 19533 5253 19567 5287
rect 21097 5253 21131 5287
rect 22937 5253 22971 5287
rect 25881 5253 25915 5287
rect 27905 5253 27939 5287
rect 6653 5185 6687 5219
rect 8217 5185 8251 5219
rect 9321 5185 9355 5219
rect 9597 5185 9631 5219
rect 10517 5185 10551 5219
rect 11529 5185 11563 5219
rect 13461 5185 13495 5219
rect 19809 5185 19843 5219
rect 19993 5185 20027 5219
rect 20913 5185 20947 5219
rect 22293 5185 22327 5219
rect 23029 5185 23063 5219
rect 23213 5185 23247 5219
rect 23397 5185 23431 5219
rect 25605 5185 25639 5219
rect 25697 5185 25731 5219
rect 27169 5185 27203 5219
rect 27629 5185 27663 5219
rect 27721 5185 27755 5219
rect 28549 5185 28583 5219
rect 28733 5185 28767 5219
rect 28917 5185 28951 5219
rect 29009 5185 29043 5219
rect 29561 5185 29595 5219
rect 29745 5185 29779 5219
rect 29929 5185 29963 5219
rect 30021 5185 30055 5219
rect 30481 5185 30515 5219
rect 30757 5185 30791 5219
rect 31125 5185 31159 5219
rect 10241 5117 10275 5151
rect 15853 5117 15887 5151
rect 16681 5117 16715 5151
rect 22385 5117 22419 5151
rect 23673 5117 23707 5151
rect 25881 5117 25915 5151
rect 27077 5117 27111 5151
rect 30573 5117 30607 5151
rect 31033 5117 31067 5151
rect 13277 5049 13311 5083
rect 19901 5049 19935 5083
rect 27905 5049 27939 5083
rect 29285 5049 29319 5083
rect 29837 5049 29871 5083
rect 30665 5049 30699 5083
rect 9137 4981 9171 5015
rect 11161 4981 11195 5015
rect 16405 4981 16439 5015
rect 23489 4981 23523 5015
rect 30297 4981 30331 5015
rect 9873 4777 9907 4811
rect 10964 4777 10998 4811
rect 12449 4777 12483 4811
rect 15945 4777 15979 4811
rect 16589 4777 16623 4811
rect 20177 4777 20211 4811
rect 20361 4777 20395 4811
rect 23489 4777 23523 4811
rect 24409 4777 24443 4811
rect 25697 4777 25731 4811
rect 26065 4777 26099 4811
rect 27537 4777 27571 4811
rect 29653 4777 29687 4811
rect 30021 4777 30055 4811
rect 30297 4777 30331 4811
rect 10701 4641 10735 4675
rect 14197 4641 14231 4675
rect 19533 4641 19567 4675
rect 24685 4641 24719 4675
rect 26617 4641 26651 4675
rect 27077 4641 27111 4675
rect 27997 4641 28031 4675
rect 28641 4641 28675 4675
rect 1777 4573 1811 4607
rect 10057 4573 10091 4607
rect 10241 4573 10275 4607
rect 16037 4573 16071 4607
rect 16313 4573 16347 4607
rect 16405 4573 16439 4607
rect 19441 4573 19475 4607
rect 21281 4573 21315 4607
rect 21833 4573 21867 4607
rect 23213 4573 23247 4607
rect 24593 4573 24627 4607
rect 24777 4573 24811 4607
rect 24869 4573 24903 4607
rect 25053 4573 25087 4607
rect 25145 4573 25179 4607
rect 25329 4573 25363 4607
rect 25605 4573 25639 4607
rect 26157 4573 26191 4607
rect 26341 4573 26375 4607
rect 26709 4573 26743 4607
rect 27353 4573 27387 4607
rect 27905 4573 27939 4607
rect 29561 4573 29595 4607
rect 30113 4573 30147 4607
rect 30297 4573 30331 4607
rect 1409 4505 1443 4539
rect 14473 4505 14507 4539
rect 16221 4505 16255 4539
rect 19993 4505 20027 4539
rect 20209 4505 20243 4539
rect 23305 4505 23339 4539
rect 23489 4505 23523 4539
rect 25513 4505 25547 4539
rect 26249 4505 26283 4539
rect 27169 4505 27203 4539
rect 19809 4437 19843 4471
rect 26433 4437 26467 4471
rect 9781 4233 9815 4267
rect 14565 4233 14599 4267
rect 27905 4233 27939 4267
rect 8309 4165 8343 4199
rect 8033 4097 8067 4131
rect 14381 4097 14415 4131
rect 24961 4097 24995 4131
rect 25145 4097 25179 4131
rect 25237 4097 25271 4131
rect 25421 4097 25455 4131
rect 27813 4097 27847 4131
rect 27997 4097 28031 4131
rect 25329 4029 25363 4063
rect 25145 3961 25179 3995
rect 37565 3077 37599 3111
rect 1961 3009 1995 3043
rect 2421 3009 2455 3043
rect 12541 3009 12575 3043
rect 13185 3009 13219 3043
rect 15117 3009 15151 3043
rect 17233 3009 17267 3043
rect 19993 3009 20027 3043
rect 1777 2805 1811 2839
rect 2237 2805 2271 2839
rect 12357 2805 12391 2839
rect 13001 2805 13035 2839
rect 14933 2805 14967 2839
rect 17417 2805 17451 2839
rect 19809 2805 19843 2839
rect 37657 2805 37691 2839
rect 8677 2601 8711 2635
rect 11161 2601 11195 2635
rect 37657 2533 37691 2567
rect 1777 2397 1811 2431
rect 2421 2397 2455 2431
rect 4353 2397 4387 2431
rect 6929 2397 6963 2431
rect 8493 2397 8527 2431
rect 13093 2397 13127 2431
rect 15025 2397 15059 2431
rect 17601 2397 17635 2431
rect 19809 2397 19843 2431
rect 37473 2397 37507 2431
rect 1409 2329 1443 2363
rect 2053 2329 2087 2363
rect 3985 2329 4019 2363
rect 6561 2329 6595 2363
rect 11253 2329 11287 2363
rect 19441 2329 19475 2363
rect 27077 2329 27111 2363
rect 13185 2261 13219 2295
rect 15301 2261 15335 2295
rect 17693 2261 17727 2295
rect 27169 2261 27203 2295
<< metal1 >>
rect 1104 39194 38272 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 38272 39194
rect 1104 39120 38272 39142
rect 14 39040 20 39092
rect 72 39080 78 39092
rect 1489 39083 1547 39089
rect 1489 39080 1501 39083
rect 72 39052 1501 39080
rect 72 39040 78 39052
rect 1489 39049 1501 39052
rect 1535 39049 1547 39083
rect 1489 39043 1547 39049
rect 4890 39040 4896 39092
rect 4948 39040 4954 39092
rect 9030 39040 9036 39092
rect 9088 39080 9094 39092
rect 9309 39083 9367 39089
rect 9309 39080 9321 39083
rect 9088 39052 9321 39080
rect 9088 39040 9094 39052
rect 9309 39049 9321 39052
rect 9355 39049 9367 39083
rect 9309 39043 9367 39049
rect 11054 39040 11060 39092
rect 11112 39080 11118 39092
rect 11609 39083 11667 39089
rect 11609 39080 11621 39083
rect 11112 39052 11621 39080
rect 11112 39040 11118 39052
rect 11609 39049 11621 39052
rect 11655 39049 11667 39083
rect 11609 39043 11667 39049
rect 13170 39040 13176 39092
rect 13228 39040 13234 39092
rect 17402 39040 17408 39092
rect 17460 39080 17466 39092
rect 17773 39083 17831 39089
rect 17773 39080 17785 39083
rect 17460 39052 17785 39080
rect 17460 39040 17466 39052
rect 17773 39049 17785 39052
rect 17819 39049 17831 39083
rect 17773 39043 17831 39049
rect 21910 39040 21916 39092
rect 21968 39080 21974 39092
rect 22097 39083 22155 39089
rect 22097 39080 22109 39083
rect 21968 39052 22109 39080
rect 21968 39040 21974 39052
rect 22097 39049 22109 39052
rect 22143 39049 22155 39083
rect 22097 39043 22155 39049
rect 26418 39040 26424 39092
rect 26476 39080 26482 39092
rect 27157 39083 27215 39089
rect 27157 39080 27169 39083
rect 26476 39052 27169 39080
rect 26476 39040 26482 39052
rect 27157 39049 27169 39052
rect 27203 39049 27215 39083
rect 27157 39043 27215 39049
rect 33134 39040 33140 39092
rect 33192 39040 33198 39092
rect 35434 39040 35440 39092
rect 35492 39080 35498 39092
rect 35713 39083 35771 39089
rect 35713 39080 35725 39083
rect 35492 39052 35725 39080
rect 35492 39040 35498 39052
rect 35713 39049 35725 39052
rect 35759 39049 35771 39083
rect 35713 39043 35771 39049
rect 11885 39015 11943 39021
rect 11885 38981 11897 39015
rect 11931 39012 11943 39015
rect 12342 39012 12348 39024
rect 11931 38984 12348 39012
rect 11931 38981 11943 38984
rect 11885 38975 11943 38981
rect 12342 38972 12348 38984
rect 12400 38972 12406 39024
rect 15470 38972 15476 39024
rect 15528 39012 15534 39024
rect 15749 39015 15807 39021
rect 15749 39012 15761 39015
rect 15528 38984 15761 39012
rect 15528 38972 15534 38984
rect 15749 38981 15761 38984
rect 15795 38981 15807 39015
rect 15749 38975 15807 38981
rect 30926 38972 30932 39024
rect 30984 39012 30990 39024
rect 31205 39015 31263 39021
rect 31205 39012 31217 39015
rect 30984 38984 31217 39012
rect 30984 38972 30990 38984
rect 31205 38981 31217 38984
rect 31251 38981 31263 39015
rect 31205 38975 31263 38981
rect 1762 38904 1768 38956
rect 1820 38904 1826 38956
rect 5074 38904 5080 38956
rect 5132 38904 5138 38956
rect 9214 38904 9220 38956
rect 9272 38904 9278 38956
rect 12066 38904 12072 38956
rect 12124 38904 12130 38956
rect 12434 38904 12440 38956
rect 12492 38944 12498 38956
rect 12989 38947 13047 38953
rect 12989 38944 13001 38947
rect 12492 38916 13001 38944
rect 12492 38904 12498 38916
rect 12989 38913 13001 38916
rect 13035 38913 13047 38947
rect 12989 38907 13047 38913
rect 17954 38904 17960 38956
rect 18012 38904 18018 38956
rect 19426 38904 19432 38956
rect 19484 38904 19490 38956
rect 20070 38904 20076 38956
rect 20128 38904 20134 38956
rect 22370 38904 22376 38956
rect 22428 38904 22434 38956
rect 27062 38904 27068 38956
rect 27120 38904 27126 38956
rect 27706 38904 27712 38956
rect 27764 38904 27770 38956
rect 33042 38904 33048 38956
rect 33100 38904 33106 38956
rect 35618 38904 35624 38956
rect 35676 38904 35682 38956
rect 37366 38904 37372 38956
rect 37424 38944 37430 38956
rect 37461 38947 37519 38953
rect 37461 38944 37473 38947
rect 37424 38916 37473 38944
rect 37424 38904 37430 38916
rect 37461 38913 37473 38916
rect 37507 38913 37519 38947
rect 37461 38907 37519 38913
rect 20346 38836 20352 38888
rect 20404 38836 20410 38888
rect 15562 38768 15568 38820
rect 15620 38768 15626 38820
rect 29730 38768 29736 38820
rect 29788 38808 29794 38820
rect 31021 38811 31079 38817
rect 31021 38808 31033 38811
rect 29788 38780 31033 38808
rect 29788 38768 29794 38780
rect 31021 38777 31033 38780
rect 31067 38777 31079 38811
rect 31021 38771 31079 38777
rect 37642 38768 37648 38820
rect 37700 38768 37706 38820
rect 12253 38743 12311 38749
rect 12253 38709 12265 38743
rect 12299 38740 12311 38743
rect 12802 38740 12808 38752
rect 12299 38712 12808 38740
rect 12299 38709 12311 38712
rect 12253 38703 12311 38709
rect 12802 38700 12808 38712
rect 12860 38700 12866 38752
rect 19610 38700 19616 38752
rect 19668 38700 19674 38752
rect 27614 38700 27620 38752
rect 27672 38700 27678 38752
rect 1104 38650 38272 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 38272 38650
rect 1104 38576 38272 38598
rect 4985 38539 5043 38545
rect 4985 38505 4997 38539
rect 5031 38536 5043 38539
rect 5074 38536 5080 38548
rect 5031 38508 5080 38536
rect 5031 38505 5043 38508
rect 4985 38499 5043 38505
rect 5074 38496 5080 38508
rect 5132 38496 5138 38548
rect 8757 38539 8815 38545
rect 8757 38505 8769 38539
rect 8803 38536 8815 38539
rect 9214 38536 9220 38548
rect 8803 38508 9220 38536
rect 8803 38505 8815 38508
rect 8757 38499 8815 38505
rect 9214 38496 9220 38508
rect 9272 38496 9278 38548
rect 17954 38496 17960 38548
rect 18012 38536 18018 38548
rect 18325 38539 18383 38545
rect 18325 38536 18337 38539
rect 18012 38508 18337 38536
rect 18012 38496 18018 38508
rect 18325 38505 18337 38508
rect 18371 38505 18383 38539
rect 27706 38536 27712 38548
rect 18325 38499 18383 38505
rect 18524 38508 20576 38536
rect 11057 38403 11115 38409
rect 11057 38369 11069 38403
rect 11103 38369 11115 38403
rect 11057 38363 11115 38369
rect 5166 38292 5172 38344
rect 5224 38292 5230 38344
rect 8570 38292 8576 38344
rect 8628 38292 8634 38344
rect 9030 38292 9036 38344
rect 9088 38292 9094 38344
rect 9125 38335 9183 38341
rect 9125 38301 9137 38335
rect 9171 38332 9183 38335
rect 9309 38335 9367 38341
rect 9309 38332 9321 38335
rect 9171 38304 9321 38332
rect 9171 38301 9183 38304
rect 9125 38295 9183 38301
rect 9309 38301 9321 38304
rect 9355 38301 9367 38335
rect 11072 38332 11100 38363
rect 11330 38332 11336 38344
rect 11072 38304 11336 38332
rect 9309 38295 9367 38301
rect 11330 38292 11336 38304
rect 11388 38292 11394 38344
rect 13081 38335 13139 38341
rect 13081 38301 13093 38335
rect 13127 38332 13139 38335
rect 13265 38335 13323 38341
rect 13265 38332 13277 38335
rect 13127 38304 13277 38332
rect 13127 38301 13139 38304
rect 13081 38295 13139 38301
rect 13265 38301 13277 38304
rect 13311 38301 13323 38335
rect 13265 38295 13323 38301
rect 13357 38335 13415 38341
rect 13357 38301 13369 38335
rect 13403 38332 13415 38335
rect 13722 38332 13728 38344
rect 13403 38304 13728 38332
rect 13403 38301 13415 38304
rect 13357 38295 13415 38301
rect 13722 38292 13728 38304
rect 13780 38292 13786 38344
rect 18524 38341 18552 38508
rect 19521 38403 19579 38409
rect 19521 38369 19533 38403
rect 19567 38400 19579 38403
rect 19610 38400 19616 38412
rect 19567 38372 19616 38400
rect 19567 38369 19579 38372
rect 19521 38363 19579 38369
rect 19610 38360 19616 38372
rect 19668 38360 19674 38412
rect 20548 38400 20576 38508
rect 25056 38508 27712 38536
rect 24854 38400 24860 38412
rect 20548 38372 24860 38400
rect 24854 38360 24860 38372
rect 24912 38360 24918 38412
rect 18509 38335 18567 38341
rect 18509 38301 18521 38335
rect 18555 38301 18567 38335
rect 18509 38295 18567 38301
rect 18877 38335 18935 38341
rect 18877 38301 18889 38335
rect 18923 38301 18935 38335
rect 18877 38295 18935 38301
rect 18969 38335 19027 38341
rect 18969 38301 18981 38335
rect 19015 38332 19027 38335
rect 19245 38335 19303 38341
rect 19245 38332 19257 38335
rect 19015 38304 19257 38332
rect 19015 38301 19027 38304
rect 18969 38295 19027 38301
rect 19245 38301 19257 38304
rect 19291 38301 19303 38335
rect 20806 38332 20812 38344
rect 20654 38304 20812 38332
rect 19245 38295 19303 38301
rect 9582 38224 9588 38276
rect 9640 38224 9646 38276
rect 10226 38224 10232 38276
rect 10284 38224 10290 38276
rect 11054 38224 11060 38276
rect 11112 38264 11118 38276
rect 11112 38236 11638 38264
rect 11112 38224 11118 38236
rect 12802 38224 12808 38276
rect 12860 38224 12866 38276
rect 12894 38224 12900 38276
rect 12952 38264 12958 38276
rect 18892 38264 18920 38295
rect 20806 38292 20812 38304
rect 20864 38292 20870 38344
rect 21266 38292 21272 38344
rect 21324 38292 21330 38344
rect 25056 38341 25084 38508
rect 27706 38496 27712 38508
rect 27764 38536 27770 38548
rect 32217 38539 32275 38545
rect 27764 38508 29592 38536
rect 27764 38496 27770 38508
rect 26050 38360 26056 38412
rect 26108 38400 26114 38412
rect 27249 38403 27307 38409
rect 26108 38372 27200 38400
rect 26108 38360 26114 38372
rect 21545 38335 21603 38341
rect 21545 38301 21557 38335
rect 21591 38301 21603 38335
rect 21545 38295 21603 38301
rect 21637 38335 21695 38341
rect 21637 38301 21649 38335
rect 21683 38332 21695 38335
rect 21821 38335 21879 38341
rect 21821 38332 21833 38335
rect 21683 38304 21833 38332
rect 21683 38301 21695 38304
rect 21637 38295 21695 38301
rect 21821 38301 21833 38304
rect 21867 38301 21879 38335
rect 21821 38295 21879 38301
rect 25041 38335 25099 38341
rect 25041 38301 25053 38335
rect 25087 38301 25099 38335
rect 25041 38295 25099 38301
rect 25133 38335 25191 38341
rect 25133 38301 25145 38335
rect 25179 38332 25191 38335
rect 25317 38335 25375 38341
rect 25317 38332 25329 38335
rect 25179 38304 25329 38332
rect 25179 38301 25191 38304
rect 25133 38295 25191 38301
rect 25317 38301 25329 38304
rect 25363 38301 25375 38335
rect 25317 38295 25375 38301
rect 21560 38264 21588 38295
rect 22097 38267 22155 38273
rect 22097 38264 22109 38267
rect 12952 38236 18920 38264
rect 20824 38236 21588 38264
rect 21744 38236 22109 38264
rect 12952 38224 12958 38236
rect 11333 38199 11391 38205
rect 11333 38165 11345 38199
rect 11379 38196 11391 38199
rect 11882 38196 11888 38208
rect 11379 38168 11888 38196
rect 11379 38165 11391 38168
rect 11333 38159 11391 38165
rect 11882 38156 11888 38168
rect 11940 38156 11946 38208
rect 13722 38156 13728 38208
rect 13780 38196 13786 38208
rect 20824 38196 20852 38236
rect 13780 38168 20852 38196
rect 13780 38156 13786 38168
rect 20990 38156 20996 38208
rect 21048 38156 21054 38208
rect 21453 38199 21511 38205
rect 21453 38165 21465 38199
rect 21499 38196 21511 38199
rect 21744 38196 21772 38236
rect 22097 38233 22109 38236
rect 22143 38233 22155 38267
rect 22097 38227 22155 38233
rect 22480 38236 22586 38264
rect 23492 38236 25544 38264
rect 21499 38168 21772 38196
rect 21499 38165 21511 38168
rect 21453 38159 21511 38165
rect 22002 38156 22008 38208
rect 22060 38196 22066 38208
rect 22480 38196 22508 38236
rect 23492 38196 23520 38236
rect 22060 38168 23520 38196
rect 23569 38199 23627 38205
rect 22060 38156 22066 38168
rect 23569 38165 23581 38199
rect 23615 38196 23627 38199
rect 24026 38196 24032 38208
rect 23615 38168 24032 38196
rect 23615 38165 23627 38168
rect 23569 38159 23627 38165
rect 24026 38156 24032 38168
rect 24084 38156 24090 38208
rect 25516 38196 25544 38236
rect 25590 38224 25596 38276
rect 25648 38224 25654 38276
rect 26050 38264 26056 38276
rect 25976 38236 26056 38264
rect 25976 38196 26004 38236
rect 26050 38224 26056 38236
rect 26108 38224 26114 38276
rect 25516 38168 26004 38196
rect 26970 38156 26976 38208
rect 27028 38196 27034 38208
rect 27065 38199 27123 38205
rect 27065 38196 27077 38199
rect 27028 38168 27077 38196
rect 27028 38156 27034 38168
rect 27065 38165 27077 38168
rect 27111 38165 27123 38199
rect 27172 38196 27200 38372
rect 27249 38369 27261 38403
rect 27295 38400 27307 38403
rect 27614 38400 27620 38412
rect 27295 38372 27620 38400
rect 27295 38369 27307 38372
rect 27249 38363 27307 38369
rect 27614 38360 27620 38372
rect 27672 38360 27678 38412
rect 29564 38344 29592 38508
rect 32217 38505 32229 38539
rect 32263 38536 32275 38539
rect 33042 38536 33048 38548
rect 32263 38508 33048 38536
rect 32263 38505 32275 38508
rect 32217 38499 32275 38505
rect 33042 38496 33048 38508
rect 33100 38496 33106 38548
rect 34885 38539 34943 38545
rect 34885 38505 34897 38539
rect 34931 38536 34943 38539
rect 35618 38536 35624 38548
rect 34931 38508 35624 38536
rect 34931 38505 34943 38508
rect 34885 38499 34943 38505
rect 35618 38496 35624 38508
rect 35676 38496 35682 38548
rect 37829 38539 37887 38545
rect 37829 38505 37841 38539
rect 37875 38536 37887 38539
rect 37918 38536 37924 38548
rect 37875 38508 37924 38536
rect 37875 38505 37887 38508
rect 37829 38499 37887 38505
rect 37918 38496 37924 38508
rect 37976 38496 37982 38548
rect 32674 38360 32680 38412
rect 32732 38400 32738 38412
rect 32732 38372 37596 38400
rect 32732 38360 32738 38372
rect 29546 38292 29552 38344
rect 29604 38292 29610 38344
rect 29638 38292 29644 38344
rect 29696 38292 29702 38344
rect 31662 38292 31668 38344
rect 31720 38332 31726 38344
rect 32033 38335 32091 38341
rect 32033 38332 32045 38335
rect 31720 38304 32045 38332
rect 31720 38292 31726 38304
rect 32033 38301 32045 38304
rect 32079 38301 32091 38335
rect 32033 38295 32091 38301
rect 34701 38335 34759 38341
rect 34701 38301 34713 38335
rect 34747 38301 34759 38335
rect 34701 38295 34759 38301
rect 27522 38224 27528 38276
rect 27580 38224 27586 38276
rect 27908 38236 28014 38264
rect 27908 38196 27936 38236
rect 29270 38224 29276 38276
rect 29328 38224 29334 38276
rect 29454 38224 29460 38276
rect 29512 38264 29518 38276
rect 29512 38236 31754 38264
rect 29512 38224 29518 38236
rect 28534 38196 28540 38208
rect 27172 38168 28540 38196
rect 27065 38159 27123 38165
rect 28534 38156 28540 38168
rect 28592 38196 28598 38208
rect 30374 38196 30380 38208
rect 28592 38168 30380 38196
rect 28592 38156 28598 38168
rect 30374 38156 30380 38168
rect 30432 38156 30438 38208
rect 31726 38196 31754 38236
rect 34716 38196 34744 38295
rect 37568 38273 37596 38372
rect 37553 38267 37611 38273
rect 37553 38233 37565 38267
rect 37599 38233 37611 38267
rect 37553 38227 37611 38233
rect 31726 38168 34744 38196
rect 1104 38106 38272 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 38272 38106
rect 1104 38032 38272 38054
rect 9582 37952 9588 38004
rect 9640 37992 9646 38004
rect 9769 37995 9827 38001
rect 9769 37992 9781 37995
rect 9640 37964 9781 37992
rect 9640 37952 9646 37964
rect 9769 37961 9781 37964
rect 9815 37961 9827 37995
rect 9769 37955 9827 37961
rect 10229 37995 10287 38001
rect 10229 37961 10241 37995
rect 10275 37961 10287 37995
rect 10229 37955 10287 37961
rect 9953 37859 10011 37865
rect 9953 37825 9965 37859
rect 9999 37856 10011 37859
rect 10244 37856 10272 37955
rect 12066 37952 12072 38004
rect 12124 37992 12130 38004
rect 12253 37995 12311 38001
rect 12253 37992 12265 37995
rect 12124 37964 12265 37992
rect 12124 37952 12130 37964
rect 12253 37961 12265 37964
rect 12299 37961 12311 37995
rect 12253 37955 12311 37961
rect 12342 37952 12348 38004
rect 12400 37952 12406 38004
rect 15286 37992 15292 38004
rect 13740 37964 15292 37992
rect 10686 37884 10692 37936
rect 10744 37924 10750 37936
rect 11793 37927 11851 37933
rect 11793 37924 11805 37927
rect 10744 37896 11805 37924
rect 10744 37884 10750 37896
rect 11793 37893 11805 37896
rect 11839 37893 11851 37927
rect 11793 37887 11851 37893
rect 11882 37884 11888 37936
rect 11940 37924 11946 37936
rect 11940 37896 13216 37924
rect 11940 37884 11946 37896
rect 9999 37828 10272 37856
rect 10597 37859 10655 37865
rect 9999 37825 10011 37828
rect 9953 37819 10011 37825
rect 10597 37825 10609 37859
rect 10643 37856 10655 37859
rect 11330 37856 11336 37868
rect 10643 37828 11336 37856
rect 10643 37825 10655 37828
rect 10597 37819 10655 37825
rect 11330 37816 11336 37828
rect 11388 37816 11394 37868
rect 12526 37816 12532 37868
rect 12584 37816 12590 37868
rect 10778 37748 10784 37800
rect 10836 37748 10842 37800
rect 11698 37748 11704 37800
rect 11756 37748 11762 37800
rect 13188 37720 13216 37896
rect 13262 37816 13268 37868
rect 13320 37816 13326 37868
rect 13740 37865 13768 37964
rect 15286 37952 15292 37964
rect 15344 37952 15350 38004
rect 16298 37952 16304 38004
rect 16356 37992 16362 38004
rect 16356 37964 19334 37992
rect 16356 37952 16362 37964
rect 14027 37927 14085 37933
rect 14027 37893 14039 37927
rect 14073 37924 14085 37927
rect 14274 37924 14280 37936
rect 14073 37896 14280 37924
rect 14073 37893 14085 37896
rect 14027 37887 14085 37893
rect 14274 37884 14280 37896
rect 14332 37884 14338 37936
rect 16684 37933 16712 37964
rect 14461 37927 14519 37933
rect 14461 37893 14473 37927
rect 14507 37924 14519 37927
rect 16669 37927 16727 37933
rect 14507 37896 16620 37924
rect 14507 37893 14519 37896
rect 14461 37887 14519 37893
rect 13725 37859 13783 37865
rect 13725 37825 13737 37859
rect 13771 37825 13783 37859
rect 13725 37819 13783 37825
rect 13814 37816 13820 37868
rect 13872 37816 13878 37868
rect 14366 37865 14372 37868
rect 13909 37859 13967 37865
rect 13909 37825 13921 37859
rect 13955 37856 13967 37859
rect 13955 37828 14320 37856
rect 13955 37825 13967 37828
rect 13909 37819 13967 37825
rect 13357 37791 13415 37797
rect 13357 37757 13369 37791
rect 13403 37788 13415 37791
rect 14185 37791 14243 37797
rect 14185 37788 14197 37791
rect 13403 37760 14197 37788
rect 13403 37757 13415 37760
rect 13357 37751 13415 37757
rect 14185 37757 14197 37760
rect 14231 37757 14243 37791
rect 14292 37788 14320 37828
rect 14364 37819 14372 37865
rect 14366 37816 14372 37819
rect 14424 37816 14430 37868
rect 14550 37816 14556 37868
rect 14608 37816 14614 37868
rect 14461 37791 14519 37797
rect 14461 37788 14473 37791
rect 14292 37760 14473 37788
rect 14185 37751 14243 37757
rect 14461 37757 14473 37760
rect 14507 37757 14519 37791
rect 14461 37751 14519 37757
rect 14090 37720 14096 37732
rect 13188 37692 14096 37720
rect 14090 37680 14096 37692
rect 14148 37720 14154 37732
rect 14660 37720 14688 37896
rect 14737 37859 14795 37865
rect 14737 37825 14749 37859
rect 14783 37825 14795 37859
rect 14737 37819 14795 37825
rect 15933 37859 15991 37865
rect 15933 37825 15945 37859
rect 15979 37856 15991 37859
rect 16022 37856 16028 37868
rect 15979 37828 16028 37856
rect 15979 37825 15991 37828
rect 15933 37819 15991 37825
rect 14752 37788 14780 37819
rect 16022 37816 16028 37828
rect 16080 37816 16086 37868
rect 16114 37816 16120 37868
rect 16172 37816 16178 37868
rect 16206 37816 16212 37868
rect 16264 37816 16270 37868
rect 16301 37859 16359 37865
rect 16301 37825 16313 37859
rect 16347 37856 16359 37859
rect 16482 37856 16488 37868
rect 16347 37828 16488 37856
rect 16347 37825 16359 37828
rect 16301 37819 16359 37825
rect 16482 37816 16488 37828
rect 16540 37816 16546 37868
rect 16592 37856 16620 37896
rect 16669 37893 16681 37927
rect 16715 37893 16727 37927
rect 16669 37887 16727 37893
rect 17037 37927 17095 37933
rect 17037 37893 17049 37927
rect 17083 37924 17095 37927
rect 17405 37927 17463 37933
rect 17405 37924 17417 37927
rect 17083 37896 17417 37924
rect 17083 37893 17095 37896
rect 17037 37887 17095 37893
rect 17405 37893 17417 37896
rect 17451 37893 17463 37927
rect 19306 37924 19334 37964
rect 19426 37952 19432 38004
rect 19484 37952 19490 38004
rect 19797 37995 19855 38001
rect 19797 37961 19809 37995
rect 19843 37992 19855 37995
rect 20990 37992 20996 38004
rect 19843 37964 20996 37992
rect 19843 37961 19855 37964
rect 19797 37955 19855 37961
rect 20990 37952 20996 37964
rect 21048 37952 21054 38004
rect 21266 37952 21272 38004
rect 21324 37992 21330 38004
rect 22005 37995 22063 38001
rect 22005 37992 22017 37995
rect 21324 37964 22017 37992
rect 21324 37952 21330 37964
rect 22005 37961 22017 37964
rect 22051 37961 22063 37995
rect 22005 37955 22063 37961
rect 22462 37952 22468 38004
rect 22520 37992 22526 38004
rect 22738 37992 22744 38004
rect 22520 37964 22744 37992
rect 22520 37952 22526 37964
rect 22738 37952 22744 37964
rect 22796 37952 22802 38004
rect 24854 37952 24860 38004
rect 24912 37952 24918 38004
rect 25590 37952 25596 38004
rect 25648 37992 25654 38004
rect 26237 37995 26295 38001
rect 26237 37992 26249 37995
rect 25648 37964 26249 37992
rect 25648 37952 25654 37964
rect 26237 37961 26249 37964
rect 26283 37961 26295 37995
rect 26237 37955 26295 37961
rect 26789 37995 26847 38001
rect 26789 37961 26801 37995
rect 26835 37992 26847 37995
rect 27522 37992 27528 38004
rect 26835 37964 27528 37992
rect 26835 37961 26847 37964
rect 26789 37955 26847 37961
rect 27522 37952 27528 37964
rect 27580 37952 27586 38004
rect 27893 37995 27951 38001
rect 27893 37961 27905 37995
rect 27939 37992 27951 37995
rect 29454 37992 29460 38004
rect 27939 37964 29460 37992
rect 27939 37961 27951 37964
rect 27893 37955 27951 37961
rect 29454 37952 29460 37964
rect 29512 37952 29518 38004
rect 29638 37952 29644 38004
rect 29696 37952 29702 38004
rect 23569 37927 23627 37933
rect 19306 37896 23024 37924
rect 17405 37887 17463 37893
rect 16850 37856 16856 37868
rect 16592 37828 16856 37856
rect 16850 37816 16856 37828
rect 16908 37816 16914 37868
rect 17218 37816 17224 37868
rect 17276 37816 17282 37868
rect 17497 37859 17555 37865
rect 17497 37825 17509 37859
rect 17543 37825 17555 37859
rect 17497 37819 17555 37825
rect 17589 37859 17647 37865
rect 17589 37825 17601 37859
rect 17635 37856 17647 37859
rect 17678 37856 17684 37868
rect 17635 37828 17684 37856
rect 17635 37825 17647 37828
rect 17589 37819 17647 37825
rect 17512 37788 17540 37819
rect 17678 37816 17684 37828
rect 17736 37816 17742 37868
rect 17862 37816 17868 37868
rect 17920 37856 17926 37868
rect 20349 37859 20407 37865
rect 20349 37856 20361 37859
rect 17920 37828 20361 37856
rect 17920 37816 17926 37828
rect 20349 37825 20361 37828
rect 20395 37825 20407 37859
rect 20349 37819 20407 37825
rect 20717 37859 20775 37865
rect 20717 37825 20729 37859
rect 20763 37856 20775 37859
rect 20806 37856 20812 37868
rect 20763 37828 20812 37856
rect 20763 37825 20775 37828
rect 20717 37819 20775 37825
rect 20806 37816 20812 37828
rect 20864 37856 20870 37868
rect 22002 37856 22008 37868
rect 20864 37828 22008 37856
rect 20864 37816 20870 37828
rect 22002 37816 22008 37828
rect 22060 37816 22066 37868
rect 22373 37859 22431 37865
rect 22373 37825 22385 37859
rect 22419 37856 22431 37859
rect 22419 37828 22968 37856
rect 22419 37825 22431 37828
rect 22373 37819 22431 37825
rect 19889 37791 19947 37797
rect 14752 37760 18184 37788
rect 14148 37692 14688 37720
rect 14148 37680 14154 37692
rect 12802 37612 12808 37664
rect 12860 37652 12866 37664
rect 13541 37655 13599 37661
rect 13541 37652 13553 37655
rect 12860 37624 13553 37652
rect 12860 37612 12866 37624
rect 13541 37621 13553 37624
rect 13587 37621 13599 37655
rect 13541 37615 13599 37621
rect 16482 37612 16488 37664
rect 16540 37612 16546 37664
rect 17773 37655 17831 37661
rect 17773 37621 17785 37655
rect 17819 37652 17831 37655
rect 17954 37652 17960 37664
rect 17819 37624 17960 37652
rect 17819 37621 17831 37624
rect 17773 37615 17831 37621
rect 17954 37612 17960 37624
rect 18012 37612 18018 37664
rect 18156 37652 18184 37760
rect 19889 37757 19901 37791
rect 19935 37788 19947 37791
rect 19978 37788 19984 37800
rect 19935 37760 19984 37788
rect 19935 37757 19947 37760
rect 19889 37751 19947 37757
rect 19978 37748 19984 37760
rect 20036 37748 20042 37800
rect 20073 37791 20131 37797
rect 20073 37757 20085 37791
rect 20119 37788 20131 37791
rect 20438 37788 20444 37800
rect 20119 37760 20444 37788
rect 20119 37757 20131 37760
rect 20073 37751 20131 37757
rect 20438 37748 20444 37760
rect 20496 37748 20502 37800
rect 22646 37788 22652 37800
rect 20640 37760 22652 37788
rect 19288 37680 19294 37732
rect 19346 37720 19352 37732
rect 20640 37720 20668 37760
rect 22646 37748 22652 37760
rect 22704 37748 22710 37800
rect 19346 37692 20668 37720
rect 19346 37680 19352 37692
rect 20714 37680 20720 37732
rect 20772 37720 20778 37732
rect 22462 37720 22468 37732
rect 20772 37692 22468 37720
rect 20772 37680 20778 37692
rect 22462 37680 22468 37692
rect 22520 37680 22526 37732
rect 22940 37720 22968 37828
rect 22996 37788 23024 37896
rect 23569 37893 23581 37927
rect 23615 37924 23627 37927
rect 24397 37927 24455 37933
rect 24397 37924 24409 37927
rect 23615 37896 24409 37924
rect 23615 37893 23627 37896
rect 23569 37887 23627 37893
rect 24397 37893 24409 37896
rect 24443 37893 24455 37927
rect 24397 37887 24455 37893
rect 25774 37884 25780 37936
rect 25832 37884 25838 37936
rect 29656 37924 29684 37952
rect 25976 37896 27752 37924
rect 23106 37816 23112 37868
rect 23164 37856 23170 37868
rect 23385 37859 23443 37865
rect 23385 37856 23397 37859
rect 23164 37828 23397 37856
rect 23164 37816 23170 37828
rect 23385 37825 23397 37828
rect 23431 37825 23443 37859
rect 23385 37819 23443 37825
rect 23658 37816 23664 37868
rect 23716 37816 23722 37868
rect 23750 37816 23756 37868
rect 23808 37816 23814 37868
rect 24029 37859 24087 37865
rect 24029 37825 24041 37859
rect 24075 37825 24087 37859
rect 24029 37819 24087 37825
rect 24213 37859 24271 37865
rect 24213 37825 24225 37859
rect 24259 37825 24271 37859
rect 24213 37819 24271 37825
rect 25041 37859 25099 37865
rect 25041 37825 25053 37859
rect 25087 37825 25099 37859
rect 25041 37819 25099 37825
rect 24044 37788 24072 37819
rect 22996 37760 24072 37788
rect 24228 37720 24256 37819
rect 22940 37692 24256 37720
rect 25056 37720 25084 37819
rect 25314 37816 25320 37868
rect 25372 37816 25378 37868
rect 25976 37865 26004 37896
rect 25501 37859 25559 37865
rect 25501 37825 25513 37859
rect 25547 37856 25559 37859
rect 25961 37859 26019 37865
rect 25961 37856 25973 37859
rect 25547 37828 25973 37856
rect 25547 37825 25559 37828
rect 25501 37819 25559 37825
rect 25961 37825 25973 37828
rect 26007 37825 26019 37859
rect 25961 37819 26019 37825
rect 25222 37748 25228 37800
rect 25280 37748 25286 37800
rect 25516 37720 25544 37819
rect 26418 37816 26424 37868
rect 26476 37816 26482 37868
rect 26602 37816 26608 37868
rect 26660 37816 26666 37868
rect 27724 37865 27752 37896
rect 29104 37896 29684 37924
rect 27709 37859 27767 37865
rect 27709 37825 27721 37859
rect 27755 37856 27767 37859
rect 28169 37859 28227 37865
rect 28169 37856 28181 37859
rect 27755 37828 28181 37856
rect 27755 37825 27767 37828
rect 27709 37819 27767 37825
rect 28169 37825 28181 37828
rect 28215 37825 28227 37859
rect 28169 37819 28227 37825
rect 28813 37859 28871 37865
rect 28813 37825 28825 37859
rect 28859 37856 28871 37859
rect 28994 37856 29000 37868
rect 28859 37828 29000 37856
rect 28859 37825 28871 37828
rect 28813 37819 28871 37825
rect 28994 37816 29000 37828
rect 29052 37816 29058 37868
rect 29104 37865 29132 37896
rect 30374 37884 30380 37936
rect 30432 37884 30438 37936
rect 29089 37859 29147 37865
rect 29089 37825 29101 37859
rect 29135 37825 29147 37859
rect 29089 37819 29147 37825
rect 31202 37816 31208 37868
rect 31260 37816 31266 37868
rect 25590 37748 25596 37800
rect 25648 37788 25654 37800
rect 25685 37791 25743 37797
rect 25685 37788 25697 37791
rect 25648 37760 25697 37788
rect 25648 37748 25654 37760
rect 25685 37757 25697 37760
rect 25731 37757 25743 37791
rect 25685 37751 25743 37757
rect 26142 37748 26148 37800
rect 26200 37748 26206 37800
rect 27062 37748 27068 37800
rect 27120 37788 27126 37800
rect 27525 37791 27583 37797
rect 27525 37788 27537 37791
rect 27120 37760 27537 37788
rect 27120 37748 27126 37760
rect 27525 37757 27537 37760
rect 27571 37757 27583 37791
rect 27525 37751 27583 37757
rect 27982 37748 27988 37800
rect 28040 37748 28046 37800
rect 29365 37791 29423 37797
rect 29365 37788 29377 37791
rect 29012 37760 29377 37788
rect 29012 37729 29040 37760
rect 29365 37757 29377 37760
rect 29411 37757 29423 37791
rect 29365 37751 29423 37757
rect 29454 37748 29460 37800
rect 29512 37788 29518 37800
rect 30837 37791 30895 37797
rect 30837 37788 30849 37791
rect 29512 37760 30849 37788
rect 29512 37748 29518 37760
rect 30837 37757 30849 37760
rect 30883 37757 30895 37791
rect 30837 37751 30895 37757
rect 31662 37748 31668 37800
rect 31720 37748 31726 37800
rect 28997 37723 29055 37729
rect 25056 37692 25728 37720
rect 24044 37664 24072 37692
rect 25700 37664 25728 37692
rect 28997 37689 29009 37723
rect 29043 37689 29055 37723
rect 31680 37720 31708 37748
rect 28997 37683 29055 37689
rect 30392 37692 31708 37720
rect 22370 37652 22376 37664
rect 18156 37624 22376 37652
rect 22370 37612 22376 37624
rect 22428 37612 22434 37664
rect 23934 37612 23940 37664
rect 23992 37612 23998 37664
rect 24026 37612 24032 37664
rect 24084 37612 24090 37664
rect 25682 37612 25688 37664
rect 25740 37612 25746 37664
rect 28353 37655 28411 37661
rect 28353 37621 28365 37655
rect 28399 37652 28411 37655
rect 30392 37652 30420 37692
rect 28399 37624 30420 37652
rect 28399 37621 28411 37624
rect 28353 37615 28411 37621
rect 30926 37612 30932 37664
rect 30984 37652 30990 37664
rect 31021 37655 31079 37661
rect 31021 37652 31033 37655
rect 30984 37624 31033 37652
rect 30984 37612 30990 37624
rect 31021 37621 31033 37624
rect 31067 37621 31079 37655
rect 31021 37615 31079 37621
rect 1104 37562 38272 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38272 37562
rect 1104 37488 38272 37510
rect 9582 37408 9588 37460
rect 9640 37448 9646 37460
rect 11054 37448 11060 37460
rect 9640 37420 11060 37448
rect 9640 37408 9646 37420
rect 11054 37408 11060 37420
rect 11112 37408 11118 37460
rect 16482 37408 16488 37460
rect 16540 37448 16546 37460
rect 17773 37451 17831 37457
rect 17773 37448 17785 37451
rect 16540 37420 17785 37448
rect 16540 37408 16546 37420
rect 17773 37417 17785 37420
rect 17819 37417 17831 37451
rect 17773 37411 17831 37417
rect 17862 37408 17868 37460
rect 17920 37408 17926 37460
rect 22370 37408 22376 37460
rect 22428 37448 22434 37460
rect 26053 37451 26111 37457
rect 22428 37420 26004 37448
rect 22428 37408 22434 37420
rect 17880 37380 17908 37408
rect 24854 37380 24860 37392
rect 12406 37352 17908 37380
rect 22848 37352 24860 37380
rect 1673 37315 1731 37321
rect 1673 37281 1685 37315
rect 1719 37312 1731 37315
rect 9582 37312 9588 37324
rect 1719 37284 9588 37312
rect 1719 37281 1731 37284
rect 1673 37275 1731 37281
rect 9582 37272 9588 37284
rect 9640 37312 9646 37324
rect 12406 37312 12434 37352
rect 9640 37284 12434 37312
rect 9640 37272 9646 37284
rect 15838 37272 15844 37324
rect 15896 37312 15902 37324
rect 16022 37312 16028 37324
rect 15896 37284 16028 37312
rect 15896 37272 15902 37284
rect 16022 37272 16028 37284
rect 16080 37312 16086 37324
rect 16080 37284 17816 37312
rect 16080 37272 16086 37284
rect 8294 37204 8300 37256
rect 8352 37204 8358 37256
rect 8573 37247 8631 37253
rect 8573 37213 8585 37247
rect 8619 37213 8631 37247
rect 8573 37207 8631 37213
rect 8665 37247 8723 37253
rect 8665 37213 8677 37247
rect 8711 37244 8723 37247
rect 8941 37247 8999 37253
rect 8941 37244 8953 37247
rect 8711 37216 8953 37244
rect 8711 37213 8723 37216
rect 8665 37207 8723 37213
rect 8941 37213 8953 37216
rect 8987 37213 8999 37247
rect 8941 37207 8999 37213
rect 934 37136 940 37188
rect 992 37176 998 37188
rect 1489 37179 1547 37185
rect 1489 37176 1501 37179
rect 992 37148 1501 37176
rect 992 37136 998 37148
rect 1489 37145 1501 37148
rect 1535 37145 1547 37179
rect 1489 37139 1547 37145
rect 7190 37136 7196 37188
rect 7248 37176 7254 37188
rect 8588 37176 8616 37207
rect 10226 37204 10232 37256
rect 10284 37244 10290 37256
rect 17788 37244 17816 37284
rect 17862 37272 17868 37324
rect 17920 37272 17926 37324
rect 22848 37312 22876 37352
rect 24854 37340 24860 37352
rect 24912 37340 24918 37392
rect 25976 37380 26004 37420
rect 26053 37417 26065 37451
rect 26099 37448 26111 37451
rect 26418 37448 26424 37460
rect 26099 37420 26424 37448
rect 26099 37417 26111 37420
rect 26053 37411 26111 37417
rect 26418 37408 26424 37420
rect 26476 37408 26482 37460
rect 26602 37408 26608 37460
rect 26660 37448 26666 37460
rect 27341 37451 27399 37457
rect 27341 37448 27353 37451
rect 26660 37420 27353 37448
rect 26660 37408 26666 37420
rect 27341 37417 27353 37420
rect 27387 37417 27399 37451
rect 27341 37411 27399 37417
rect 25976 37352 26556 37380
rect 17972 37284 22876 37312
rect 17972 37244 18000 37284
rect 22922 37272 22928 37324
rect 22980 37272 22986 37324
rect 23474 37272 23480 37324
rect 23532 37272 23538 37324
rect 10284 37216 10350 37244
rect 17788 37216 18000 37244
rect 18049 37247 18107 37253
rect 10284 37204 10290 37216
rect 18049 37213 18061 37247
rect 18095 37244 18107 37247
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18095 37216 18337 37244
rect 18095 37213 18107 37216
rect 18049 37207 18107 37213
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 18414 37204 18420 37256
rect 18472 37244 18478 37256
rect 18509 37247 18567 37253
rect 18509 37244 18521 37247
rect 18472 37216 18521 37244
rect 18472 37204 18478 37216
rect 18509 37213 18521 37216
rect 18555 37213 18567 37247
rect 18509 37207 18567 37213
rect 18601 37247 18659 37253
rect 18601 37213 18613 37247
rect 18647 37213 18659 37247
rect 18601 37207 18659 37213
rect 7248 37148 8616 37176
rect 9217 37179 9275 37185
rect 7248 37136 7254 37148
rect 9217 37145 9229 37179
rect 9263 37145 9275 37179
rect 9217 37139 9275 37145
rect 8481 37111 8539 37117
rect 8481 37077 8493 37111
rect 8527 37108 8539 37111
rect 9232 37108 9260 37139
rect 17770 37136 17776 37188
rect 17828 37136 17834 37188
rect 18616 37176 18644 37207
rect 20162 37204 20168 37256
rect 20220 37204 20226 37256
rect 20257 37247 20315 37253
rect 20257 37213 20269 37247
rect 20303 37244 20315 37247
rect 20441 37247 20499 37253
rect 20441 37244 20453 37247
rect 20303 37216 20453 37244
rect 20303 37213 20315 37216
rect 20257 37207 20315 37213
rect 20441 37213 20453 37216
rect 20487 37213 20499 37247
rect 20441 37207 20499 37213
rect 22738 37204 22744 37256
rect 22796 37204 22802 37256
rect 23290 37204 23296 37256
rect 23348 37204 23354 37256
rect 23492 37244 23520 37272
rect 23661 37247 23719 37253
rect 23661 37244 23673 37247
rect 23492 37216 23673 37244
rect 23661 37213 23673 37216
rect 23707 37244 23719 37247
rect 24394 37244 24400 37256
rect 23707 37216 24400 37244
rect 23707 37213 23719 37216
rect 23661 37207 23719 37213
rect 24394 37204 24400 37216
rect 24452 37204 24458 37256
rect 24872 37244 24900 37340
rect 26421 37247 26479 37253
rect 26421 37244 26433 37247
rect 24872 37216 26433 37244
rect 26421 37213 26433 37216
rect 26467 37213 26479 37247
rect 26528 37244 26556 37352
rect 26697 37315 26755 37321
rect 26697 37281 26709 37315
rect 26743 37312 26755 37315
rect 27890 37312 27896 37324
rect 26743 37284 27896 37312
rect 26743 37281 26755 37284
rect 26697 37275 26755 37281
rect 27890 37272 27896 37284
rect 27948 37272 27954 37324
rect 27985 37315 28043 37321
rect 27985 37281 27997 37315
rect 28031 37312 28043 37315
rect 28626 37312 28632 37324
rect 28031 37284 28632 37312
rect 28031 37281 28043 37284
rect 27985 37275 28043 37281
rect 28626 37272 28632 37284
rect 28684 37272 28690 37324
rect 29546 37272 29552 37324
rect 29604 37312 29610 37324
rect 30193 37315 30251 37321
rect 29604 37284 29684 37312
rect 29604 37272 29610 37284
rect 27338 37244 27344 37256
rect 26528 37216 27344 37244
rect 26421 37207 26479 37213
rect 18161 37148 18644 37176
rect 8527 37080 9260 37108
rect 8527 37077 8539 37080
rect 8481 37071 8539 37077
rect 10594 37068 10600 37120
rect 10652 37108 10658 37120
rect 10689 37111 10747 37117
rect 10689 37108 10701 37111
rect 10652 37080 10701 37108
rect 10652 37068 10658 37080
rect 10689 37077 10701 37080
rect 10735 37077 10747 37111
rect 10689 37071 10747 37077
rect 17126 37068 17132 37120
rect 17184 37108 17190 37120
rect 18161 37108 18189 37148
rect 20714 37136 20720 37188
rect 20772 37136 20778 37188
rect 22002 37176 22008 37188
rect 21942 37148 22008 37176
rect 22002 37136 22008 37148
rect 22060 37136 22066 37188
rect 22830 37176 22836 37188
rect 22204 37148 22836 37176
rect 17184 37080 18189 37108
rect 18233 37111 18291 37117
rect 17184 37068 17190 37080
rect 18233 37077 18245 37111
rect 18279 37108 18291 37111
rect 18506 37108 18512 37120
rect 18279 37080 18512 37108
rect 18279 37077 18291 37080
rect 18233 37071 18291 37077
rect 18506 37068 18512 37080
rect 18564 37068 18570 37120
rect 22204 37117 22232 37148
rect 22830 37136 22836 37148
rect 22888 37136 22894 37188
rect 23477 37179 23535 37185
rect 23477 37176 23489 37179
rect 23400 37148 23489 37176
rect 22189 37111 22247 37117
rect 22189 37077 22201 37111
rect 22235 37077 22247 37111
rect 22189 37071 22247 37077
rect 22370 37068 22376 37120
rect 22428 37068 22434 37120
rect 23400 37108 23428 37148
rect 23477 37145 23489 37148
rect 23523 37145 23535 37179
rect 23477 37139 23535 37145
rect 23566 37136 23572 37188
rect 23624 37136 23630 37188
rect 24670 37176 24676 37188
rect 23676 37148 24676 37176
rect 23676 37108 23704 37148
rect 24670 37136 24676 37148
rect 24728 37136 24734 37188
rect 26436 37176 26464 37207
rect 27338 37204 27344 37216
rect 27396 37244 27402 37256
rect 27801 37247 27859 37253
rect 27801 37244 27813 37247
rect 27396 37216 27813 37244
rect 27396 37204 27402 37216
rect 27801 37213 27813 37216
rect 27847 37244 27859 37247
rect 29270 37244 29276 37256
rect 27847 37216 29276 37244
rect 27847 37213 27859 37216
rect 27801 37207 27859 37213
rect 29270 37204 29276 37216
rect 29328 37204 29334 37256
rect 29656 37253 29684 37284
rect 30193 37281 30205 37315
rect 30239 37312 30251 37315
rect 30926 37312 30932 37324
rect 30239 37284 30932 37312
rect 30239 37281 30251 37284
rect 30193 37275 30251 37281
rect 30926 37272 30932 37284
rect 30984 37272 30990 37324
rect 29641 37247 29699 37253
rect 29641 37213 29653 37247
rect 29687 37213 29699 37247
rect 29641 37207 29699 37213
rect 29733 37247 29791 37253
rect 29733 37213 29745 37247
rect 29779 37244 29791 37247
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 29779 37216 29929 37244
rect 29779 37213 29791 37216
rect 29733 37207 29791 37213
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 29917 37207 29975 37213
rect 32582 37204 32588 37256
rect 32640 37204 32646 37256
rect 37645 37247 37703 37253
rect 37645 37213 37657 37247
rect 37691 37213 37703 37247
rect 37645 37207 37703 37213
rect 26970 37176 26976 37188
rect 26436 37148 26976 37176
rect 26970 37136 26976 37148
rect 27028 37176 27034 37188
rect 27982 37176 27988 37188
rect 27028 37148 27988 37176
rect 27028 37136 27034 37148
rect 27982 37136 27988 37148
rect 28040 37136 28046 37188
rect 30466 37136 30472 37188
rect 30524 37176 30530 37188
rect 30524 37148 30682 37176
rect 30524 37136 30530 37148
rect 31478 37136 31484 37188
rect 31536 37176 31542 37188
rect 37660 37176 37688 37207
rect 31536 37148 37688 37176
rect 31536 37136 31542 37148
rect 23400 37080 23704 37108
rect 23845 37111 23903 37117
rect 23845 37077 23857 37111
rect 23891 37108 23903 37111
rect 24578 37108 24584 37120
rect 23891 37080 24584 37108
rect 23891 37077 23903 37080
rect 23845 37071 23903 37077
rect 24578 37068 24584 37080
rect 24636 37068 24642 37120
rect 26513 37111 26571 37117
rect 26513 37077 26525 37111
rect 26559 37108 26571 37111
rect 27614 37108 27620 37120
rect 26559 37080 27620 37108
rect 26559 37077 26571 37080
rect 26513 37071 26571 37077
rect 27614 37068 27620 37080
rect 27672 37108 27678 37120
rect 27709 37111 27767 37117
rect 27709 37108 27721 37111
rect 27672 37080 27721 37108
rect 27672 37068 27678 37080
rect 27709 37077 27721 37080
rect 27755 37077 27767 37111
rect 27709 37071 27767 37077
rect 30006 37068 30012 37120
rect 30064 37108 30070 37120
rect 31665 37111 31723 37117
rect 31665 37108 31677 37111
rect 30064 37080 31677 37108
rect 30064 37068 30070 37080
rect 31665 37077 31677 37080
rect 31711 37077 31723 37111
rect 31665 37071 31723 37077
rect 32490 37068 32496 37120
rect 32548 37068 32554 37120
rect 37826 37068 37832 37120
rect 37884 37068 37890 37120
rect 1104 37018 38272 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38272 37018
rect 1104 36944 38272 36966
rect 8294 36864 8300 36916
rect 8352 36904 8358 36916
rect 9309 36907 9367 36913
rect 9309 36904 9321 36907
rect 8352 36876 9321 36904
rect 8352 36864 8358 36876
rect 9309 36873 9321 36876
rect 9355 36873 9367 36907
rect 9309 36867 9367 36873
rect 9677 36907 9735 36913
rect 9677 36873 9689 36907
rect 9723 36904 9735 36907
rect 10686 36904 10692 36916
rect 9723 36876 10692 36904
rect 9723 36873 9735 36876
rect 9677 36867 9735 36873
rect 10686 36864 10692 36876
rect 10744 36864 10750 36916
rect 20714 36864 20720 36916
rect 20772 36904 20778 36916
rect 20901 36907 20959 36913
rect 20901 36904 20913 36907
rect 20772 36876 20913 36904
rect 20772 36864 20778 36876
rect 20901 36873 20913 36876
rect 20947 36873 20959 36907
rect 22370 36904 22376 36916
rect 20901 36867 20959 36873
rect 22066 36876 22376 36904
rect 8757 36839 8815 36845
rect 8757 36805 8769 36839
rect 8803 36836 8815 36839
rect 9582 36836 9588 36848
rect 8803 36808 9588 36836
rect 8803 36805 8815 36808
rect 8757 36799 8815 36805
rect 9582 36796 9588 36808
rect 9640 36796 9646 36848
rect 9769 36839 9827 36845
rect 9769 36805 9781 36839
rect 9815 36836 9827 36839
rect 10594 36836 10600 36848
rect 9815 36808 10600 36836
rect 9815 36805 9827 36808
rect 9769 36799 9827 36805
rect 10594 36796 10600 36808
rect 10652 36796 10658 36848
rect 7285 36771 7343 36777
rect 7285 36737 7297 36771
rect 7331 36768 7343 36771
rect 7331 36740 8064 36768
rect 7331 36737 7343 36740
rect 7285 36731 7343 36737
rect 8036 36709 8064 36740
rect 14274 36728 14280 36780
rect 14332 36768 14338 36780
rect 14826 36768 14832 36780
rect 14332 36740 14832 36768
rect 14332 36728 14338 36740
rect 14826 36728 14832 36740
rect 14884 36728 14890 36780
rect 17494 36728 17500 36780
rect 17552 36768 17558 36780
rect 18414 36768 18420 36780
rect 17552 36740 18420 36768
rect 17552 36728 17558 36740
rect 18414 36728 18420 36740
rect 18472 36768 18478 36780
rect 19978 36768 19984 36780
rect 18472 36740 19984 36768
rect 18472 36728 18478 36740
rect 19978 36728 19984 36740
rect 20036 36728 20042 36780
rect 21085 36771 21143 36777
rect 21085 36737 21097 36771
rect 21131 36768 21143 36771
rect 22066 36768 22094 36876
rect 22370 36864 22376 36876
rect 22428 36864 22434 36916
rect 23584 36876 24900 36904
rect 21131 36740 22094 36768
rect 21131 36737 21143 36740
rect 21085 36731 21143 36737
rect 22462 36728 22468 36780
rect 22520 36768 22526 36780
rect 23474 36768 23480 36780
rect 22520 36740 23480 36768
rect 22520 36728 22526 36740
rect 23474 36728 23480 36740
rect 23532 36728 23538 36780
rect 8021 36703 8079 36709
rect 8021 36669 8033 36703
rect 8067 36700 8079 36703
rect 9490 36700 9496 36712
rect 8067 36672 9496 36700
rect 8067 36669 8079 36672
rect 8021 36663 8079 36669
rect 9490 36660 9496 36672
rect 9548 36660 9554 36712
rect 9858 36660 9864 36712
rect 9916 36660 9922 36712
rect 17034 36660 17040 36712
rect 17092 36700 17098 36712
rect 19150 36700 19156 36712
rect 17092 36672 19156 36700
rect 17092 36660 17098 36672
rect 19150 36660 19156 36672
rect 19208 36660 19214 36712
rect 20714 36660 20720 36712
rect 20772 36700 20778 36712
rect 23584 36700 23612 36876
rect 24029 36839 24087 36845
rect 24029 36805 24041 36839
rect 24075 36836 24087 36839
rect 24872 36836 24900 36876
rect 25130 36864 25136 36916
rect 25188 36904 25194 36916
rect 27798 36904 27804 36916
rect 25188 36876 27804 36904
rect 25188 36864 25194 36876
rect 27798 36864 27804 36876
rect 27856 36904 27862 36916
rect 28077 36907 28135 36913
rect 28077 36904 28089 36907
rect 27856 36876 28089 36904
rect 27856 36864 27862 36876
rect 28077 36873 28089 36876
rect 28123 36873 28135 36907
rect 28077 36867 28135 36873
rect 28994 36864 29000 36916
rect 29052 36904 29058 36916
rect 29181 36907 29239 36913
rect 29181 36904 29193 36907
rect 29052 36876 29193 36904
rect 29052 36864 29058 36876
rect 29181 36873 29193 36876
rect 29227 36873 29239 36907
rect 29181 36867 29239 36873
rect 30006 36864 30012 36916
rect 30064 36904 30070 36916
rect 30929 36907 30987 36913
rect 30929 36904 30941 36907
rect 30064 36876 30941 36904
rect 30064 36864 30070 36876
rect 30929 36873 30941 36876
rect 30975 36873 30987 36907
rect 30929 36867 30987 36873
rect 31202 36864 31208 36916
rect 31260 36904 31266 36916
rect 31297 36907 31355 36913
rect 31297 36904 31309 36907
rect 31260 36876 31309 36904
rect 31260 36864 31266 36876
rect 31297 36873 31309 36876
rect 31343 36873 31355 36907
rect 31297 36867 31355 36873
rect 31478 36864 31484 36916
rect 31536 36864 31542 36916
rect 32490 36864 32496 36916
rect 32548 36864 32554 36916
rect 31496 36836 31524 36864
rect 32508 36836 32536 36864
rect 24075 36808 24808 36836
rect 24872 36808 31524 36836
rect 32324 36808 32536 36836
rect 24075 36805 24087 36808
rect 24029 36799 24087 36805
rect 23845 36771 23903 36777
rect 23845 36737 23857 36771
rect 23891 36737 23903 36771
rect 23845 36731 23903 36737
rect 20772 36672 23612 36700
rect 23661 36703 23719 36709
rect 20772 36660 20778 36672
rect 23661 36669 23673 36703
rect 23707 36669 23719 36703
rect 23860 36700 23888 36731
rect 23934 36728 23940 36780
rect 23992 36768 23998 36780
rect 23992 36740 24348 36768
rect 23992 36728 23998 36740
rect 24320 36700 24348 36740
rect 24486 36728 24492 36780
rect 24544 36728 24550 36780
rect 24780 36777 24808 36808
rect 24765 36771 24823 36777
rect 24765 36737 24777 36771
rect 24811 36737 24823 36771
rect 24765 36731 24823 36737
rect 27706 36728 27712 36780
rect 27764 36728 27770 36780
rect 27985 36771 28043 36777
rect 27985 36737 27997 36771
rect 28031 36737 28043 36771
rect 27985 36731 28043 36737
rect 24581 36703 24639 36709
rect 24581 36700 24593 36703
rect 23860 36672 24164 36700
rect 24320 36672 24593 36700
rect 23661 36663 23719 36669
rect 22554 36632 22560 36644
rect 15764 36604 22560 36632
rect 15764 36576 15792 36604
rect 22554 36592 22560 36604
rect 22612 36592 22618 36644
rect 23474 36592 23480 36644
rect 23532 36632 23538 36644
rect 23676 36632 23704 36663
rect 24136 36644 24164 36672
rect 24581 36669 24593 36672
rect 24627 36669 24639 36703
rect 24581 36663 24639 36669
rect 27890 36660 27896 36712
rect 27948 36660 27954 36712
rect 28000 36700 28028 36731
rect 28258 36728 28264 36780
rect 28316 36728 28322 36780
rect 29362 36728 29368 36780
rect 29420 36768 29426 36780
rect 32324 36777 32352 36808
rect 29549 36771 29607 36777
rect 29549 36768 29561 36771
rect 29420 36740 29561 36768
rect 29420 36728 29426 36740
rect 29549 36737 29561 36740
rect 29595 36768 29607 36771
rect 30837 36771 30895 36777
rect 30837 36768 30849 36771
rect 29595 36740 30849 36768
rect 29595 36737 29607 36740
rect 29549 36731 29607 36737
rect 30837 36737 30849 36740
rect 30883 36737 30895 36771
rect 30837 36731 30895 36737
rect 32309 36771 32367 36777
rect 32309 36737 32321 36771
rect 32355 36737 32367 36771
rect 32309 36731 32367 36737
rect 28166 36700 28172 36712
rect 28000 36672 28172 36700
rect 28166 36660 28172 36672
rect 28224 36660 28230 36712
rect 29454 36660 29460 36712
rect 29512 36700 29518 36712
rect 29638 36700 29644 36712
rect 29512 36672 29644 36700
rect 29512 36660 29518 36672
rect 29638 36660 29644 36672
rect 29696 36660 29702 36712
rect 29733 36703 29791 36709
rect 29733 36669 29745 36703
rect 29779 36669 29791 36703
rect 29733 36663 29791 36669
rect 23532 36604 23704 36632
rect 23532 36592 23538 36604
rect 23934 36592 23940 36644
rect 23992 36632 23998 36644
rect 24118 36632 24124 36644
rect 23992 36604 24124 36632
rect 23992 36592 23998 36604
rect 24118 36592 24124 36604
rect 24176 36592 24182 36644
rect 25130 36632 25136 36644
rect 24504 36604 25136 36632
rect 7466 36524 7472 36576
rect 7524 36564 7530 36576
rect 7561 36567 7619 36573
rect 7561 36564 7573 36567
rect 7524 36536 7573 36564
rect 7524 36524 7530 36536
rect 7561 36533 7573 36536
rect 7607 36533 7619 36567
rect 7561 36527 7619 36533
rect 11514 36524 11520 36576
rect 11572 36564 11578 36576
rect 15654 36564 15660 36576
rect 11572 36536 15660 36564
rect 11572 36524 11578 36536
rect 15654 36524 15660 36536
rect 15712 36524 15718 36576
rect 15746 36524 15752 36576
rect 15804 36524 15810 36576
rect 17954 36524 17960 36576
rect 18012 36564 18018 36576
rect 24504 36564 24532 36604
rect 25130 36592 25136 36604
rect 25188 36592 25194 36644
rect 27908 36632 27936 36660
rect 29270 36632 29276 36644
rect 27908 36604 29276 36632
rect 29270 36592 29276 36604
rect 29328 36592 29334 36644
rect 18012 36536 24532 36564
rect 18012 36524 18018 36536
rect 24578 36524 24584 36576
rect 24636 36524 24642 36576
rect 24949 36567 25007 36573
rect 24949 36533 24961 36567
rect 24995 36564 25007 36567
rect 26234 36564 26240 36576
rect 24995 36536 26240 36564
rect 24995 36533 25007 36536
rect 24949 36527 25007 36533
rect 26234 36524 26240 36536
rect 26292 36524 26298 36576
rect 27430 36524 27436 36576
rect 27488 36564 27494 36576
rect 27617 36567 27675 36573
rect 27617 36564 27629 36567
rect 27488 36536 27629 36564
rect 27488 36524 27494 36536
rect 27617 36533 27629 36536
rect 27663 36533 27675 36567
rect 27617 36527 27675 36533
rect 28442 36524 28448 36576
rect 28500 36524 28506 36576
rect 28626 36524 28632 36576
rect 28684 36564 28690 36576
rect 29749 36564 29777 36663
rect 30650 36660 30656 36712
rect 30708 36660 30714 36712
rect 28684 36536 29777 36564
rect 30852 36564 30880 36731
rect 33686 36728 33692 36780
rect 33744 36728 33750 36780
rect 32214 36660 32220 36712
rect 32272 36700 32278 36712
rect 32585 36703 32643 36709
rect 32585 36700 32597 36703
rect 32272 36672 32597 36700
rect 32272 36660 32278 36672
rect 32585 36669 32597 36672
rect 32631 36669 32643 36703
rect 32585 36663 32643 36669
rect 33134 36564 33140 36576
rect 30852 36536 33140 36564
rect 28684 36524 28690 36536
rect 33134 36524 33140 36536
rect 33192 36524 33198 36576
rect 34054 36524 34060 36576
rect 34112 36524 34118 36576
rect 1104 36474 38272 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38272 36474
rect 1104 36400 38272 36422
rect 11793 36363 11851 36369
rect 11793 36329 11805 36363
rect 11839 36360 11851 36363
rect 12529 36363 12587 36369
rect 12529 36360 12541 36363
rect 11839 36332 12541 36360
rect 11839 36329 11851 36332
rect 11793 36323 11851 36329
rect 12529 36329 12541 36332
rect 12575 36329 12587 36363
rect 12529 36323 12587 36329
rect 13170 36320 13176 36372
rect 13228 36360 13234 36372
rect 13630 36360 13636 36372
rect 13228 36332 13636 36360
rect 13228 36320 13234 36332
rect 13630 36320 13636 36332
rect 13688 36320 13694 36372
rect 13814 36320 13820 36372
rect 13872 36360 13878 36372
rect 14277 36363 14335 36369
rect 14277 36360 14289 36363
rect 13872 36332 14289 36360
rect 13872 36320 13878 36332
rect 14277 36329 14289 36332
rect 14323 36329 14335 36363
rect 14277 36323 14335 36329
rect 14550 36320 14556 36372
rect 14608 36360 14614 36372
rect 15194 36360 15200 36372
rect 14608 36332 15200 36360
rect 14608 36320 14614 36332
rect 15194 36320 15200 36332
rect 15252 36320 15258 36372
rect 15286 36320 15292 36372
rect 15344 36320 15350 36372
rect 16485 36363 16543 36369
rect 16485 36329 16497 36363
rect 16531 36360 16543 36363
rect 16758 36360 16764 36372
rect 16531 36332 16764 36360
rect 16531 36329 16543 36332
rect 16485 36323 16543 36329
rect 16758 36320 16764 36332
rect 16816 36320 16822 36372
rect 17770 36320 17776 36372
rect 17828 36360 17834 36372
rect 18049 36363 18107 36369
rect 18049 36360 18061 36363
rect 17828 36332 18061 36360
rect 17828 36320 17834 36332
rect 18049 36329 18061 36332
rect 18095 36329 18107 36363
rect 22462 36360 22468 36372
rect 18049 36323 18107 36329
rect 18708 36332 22468 36360
rect 11698 36252 11704 36304
rect 11756 36292 11762 36304
rect 11977 36295 12035 36301
rect 11977 36292 11989 36295
rect 11756 36264 11989 36292
rect 11756 36252 11762 36264
rect 11977 36261 11989 36264
rect 12023 36261 12035 36295
rect 11977 36255 12035 36261
rect 12713 36295 12771 36301
rect 12713 36261 12725 36295
rect 12759 36261 12771 36295
rect 17126 36292 17132 36304
rect 12713 36255 12771 36261
rect 13004 36264 17132 36292
rect 6822 36184 6828 36236
rect 6880 36224 6886 36236
rect 7466 36224 7472 36236
rect 6880 36196 7472 36224
rect 6880 36184 6886 36196
rect 7466 36184 7472 36196
rect 7524 36184 7530 36236
rect 12621 36227 12679 36233
rect 10612 36196 11468 36224
rect 5718 36116 5724 36168
rect 5776 36116 5782 36168
rect 5813 36159 5871 36165
rect 5813 36125 5825 36159
rect 5859 36156 5871 36159
rect 5997 36159 6055 36165
rect 5997 36156 6009 36159
rect 5859 36128 6009 36156
rect 5859 36125 5871 36128
rect 5813 36119 5871 36125
rect 5997 36125 6009 36128
rect 6043 36125 6055 36159
rect 5997 36119 6055 36125
rect 6270 36048 6276 36100
rect 6328 36048 6334 36100
rect 7484 36088 7512 36184
rect 10612 36168 10640 36196
rect 9030 36116 9036 36168
rect 9088 36156 9094 36168
rect 9493 36159 9551 36165
rect 9493 36156 9505 36159
rect 9088 36128 9505 36156
rect 9088 36116 9094 36128
rect 9493 36125 9505 36128
rect 9539 36125 9551 36159
rect 9493 36119 9551 36125
rect 9766 36116 9772 36168
rect 9824 36116 9830 36168
rect 10226 36116 10232 36168
rect 10284 36116 10290 36168
rect 10594 36116 10600 36168
rect 10652 36116 10658 36168
rect 11241 36159 11299 36165
rect 11241 36125 11253 36159
rect 11287 36156 11299 36159
rect 11330 36156 11336 36168
rect 11287 36128 11336 36156
rect 11287 36125 11299 36128
rect 11241 36119 11299 36125
rect 11330 36116 11336 36128
rect 11388 36116 11394 36168
rect 11440 36156 11468 36196
rect 12621 36193 12633 36227
rect 12667 36224 12679 36227
rect 12728 36224 12756 36255
rect 12667 36196 12756 36224
rect 12667 36193 12679 36196
rect 12621 36187 12679 36193
rect 11514 36156 11520 36168
rect 11440 36128 11520 36156
rect 11514 36116 11520 36128
rect 11572 36116 11578 36168
rect 11609 36159 11667 36165
rect 11609 36125 11621 36159
rect 11655 36156 11667 36159
rect 11882 36156 11888 36168
rect 11655 36128 11888 36156
rect 11655 36125 11667 36128
rect 11609 36119 11667 36125
rect 11882 36116 11888 36128
rect 11940 36116 11946 36168
rect 12099 36159 12157 36165
rect 12099 36156 12111 36159
rect 12083 36125 12111 36156
rect 12145 36125 12157 36159
rect 12083 36119 12157 36125
rect 10244 36088 10272 36116
rect 7484 36074 10272 36088
rect 7498 36060 10272 36074
rect 11425 36091 11483 36097
rect 11425 36057 11437 36091
rect 11471 36057 11483 36091
rect 11425 36051 11483 36057
rect 7742 35980 7748 36032
rect 7800 35980 7806 36032
rect 9398 35980 9404 36032
rect 9456 35980 9462 36032
rect 9582 35980 9588 36032
rect 9640 35980 9646 36032
rect 11440 36020 11468 36051
rect 11790 36048 11796 36100
rect 11848 36088 11854 36100
rect 12083 36088 12111 36119
rect 12250 36116 12256 36168
rect 12308 36156 12314 36168
rect 12851 36159 12909 36165
rect 12851 36156 12863 36159
rect 12308 36128 12863 36156
rect 12308 36116 12314 36128
rect 12851 36125 12863 36128
rect 12897 36125 12909 36159
rect 12851 36119 12909 36125
rect 13004 36100 13032 36264
rect 13279 36196 14136 36224
rect 13170 36156 13176 36168
rect 13096 36128 13176 36156
rect 11848 36060 12940 36088
rect 11848 36048 11854 36060
rect 11974 36020 11980 36032
rect 11440 35992 11980 36020
rect 11974 35980 11980 35992
rect 12032 35980 12038 36032
rect 12161 36023 12219 36029
rect 12161 35989 12173 36023
rect 12207 36020 12219 36023
rect 12802 36020 12808 36032
rect 12207 35992 12808 36020
rect 12207 35989 12219 35992
rect 12161 35983 12219 35989
rect 12802 35980 12808 35992
rect 12860 35980 12866 36032
rect 12912 36020 12940 36060
rect 12986 36048 12992 36100
rect 13044 36048 13050 36100
rect 13096 36097 13124 36128
rect 13170 36116 13176 36128
rect 13228 36116 13234 36168
rect 13279 36165 13307 36196
rect 14108 36168 14136 36196
rect 13264 36159 13322 36165
rect 13264 36125 13276 36159
rect 13310 36125 13322 36159
rect 13264 36119 13322 36125
rect 13357 36159 13415 36165
rect 13357 36125 13369 36159
rect 13403 36125 13415 36159
rect 13357 36119 13415 36125
rect 13081 36091 13139 36097
rect 13081 36057 13093 36091
rect 13127 36057 13139 36091
rect 13081 36051 13139 36057
rect 13372 36020 13400 36119
rect 14090 36116 14096 36168
rect 14148 36116 14154 36168
rect 14274 36116 14280 36168
rect 14332 36116 14338 36168
rect 14369 36159 14427 36165
rect 14369 36125 14381 36159
rect 14415 36125 14427 36159
rect 14568 36156 14596 36264
rect 17126 36252 17132 36264
rect 17184 36252 17190 36304
rect 17954 36224 17960 36236
rect 15580 36196 17960 36224
rect 14645 36159 14703 36165
rect 14645 36156 14657 36159
rect 14568 36128 14657 36156
rect 14369 36119 14427 36125
rect 14645 36125 14657 36128
rect 14691 36125 14703 36159
rect 14645 36119 14703 36125
rect 14737 36159 14795 36165
rect 14737 36125 14749 36159
rect 14783 36125 14795 36159
rect 14737 36119 14795 36125
rect 12912 35992 13400 36020
rect 14384 36020 14412 36119
rect 14550 36048 14556 36100
rect 14608 36048 14614 36100
rect 14752 36088 14780 36119
rect 14826 36116 14832 36168
rect 14884 36156 14890 36168
rect 15289 36159 15347 36165
rect 15289 36156 15301 36159
rect 14884 36128 15301 36156
rect 14884 36116 14890 36128
rect 15289 36125 15301 36128
rect 15335 36125 15347 36159
rect 15289 36119 15347 36125
rect 15381 36159 15439 36165
rect 15381 36125 15393 36159
rect 15427 36156 15439 36159
rect 15580 36156 15608 36196
rect 15427 36128 15608 36156
rect 15427 36125 15439 36128
rect 15381 36119 15439 36125
rect 15654 36116 15660 36168
rect 15712 36116 15718 36168
rect 15746 36116 15752 36168
rect 15804 36116 15810 36168
rect 15933 36159 15991 36165
rect 15933 36125 15945 36159
rect 15979 36125 15991 36159
rect 15933 36119 15991 36125
rect 15102 36088 15108 36100
rect 14752 36060 15108 36088
rect 15102 36048 15108 36060
rect 15160 36048 15166 36100
rect 15562 36048 15568 36100
rect 15620 36048 15626 36100
rect 15672 36088 15700 36116
rect 15948 36088 15976 36119
rect 16206 36116 16212 36168
rect 16264 36116 16270 36168
rect 16301 36159 16359 36165
rect 16301 36125 16313 36159
rect 16347 36156 16359 36159
rect 16666 36156 16672 36168
rect 16347 36128 16672 36156
rect 16347 36125 16359 36128
rect 16301 36119 16359 36125
rect 16666 36116 16672 36128
rect 16724 36116 16730 36168
rect 16758 36116 16764 36168
rect 16816 36116 16822 36168
rect 16850 36116 16856 36168
rect 16908 36116 16914 36168
rect 17218 36116 17224 36168
rect 17276 36165 17282 36168
rect 17788 36165 17816 36196
rect 17954 36184 17960 36196
rect 18012 36184 18018 36236
rect 17276 36156 17284 36165
rect 17497 36159 17555 36165
rect 17276 36128 17321 36156
rect 17276 36119 17284 36128
rect 17497 36125 17509 36159
rect 17543 36125 17555 36159
rect 17497 36119 17555 36125
rect 17773 36159 17831 36165
rect 17773 36125 17785 36159
rect 17819 36125 17831 36159
rect 17773 36119 17831 36125
rect 17276 36116 17282 36119
rect 15672 36060 15976 36088
rect 15838 36020 15844 36032
rect 14384 35992 15844 36020
rect 15838 35980 15844 35992
rect 15896 35980 15902 36032
rect 15948 36020 15976 36060
rect 16114 36048 16120 36100
rect 16172 36048 16178 36100
rect 17034 36048 17040 36100
rect 17092 36048 17098 36100
rect 17126 36048 17132 36100
rect 17184 36048 17190 36100
rect 17512 36088 17540 36119
rect 17862 36116 17868 36168
rect 17920 36116 17926 36168
rect 18046 36116 18052 36168
rect 18104 36156 18110 36168
rect 18708 36165 18736 36332
rect 22462 36320 22468 36332
rect 22520 36320 22526 36372
rect 23014 36320 23020 36372
rect 23072 36360 23078 36372
rect 23566 36360 23572 36372
rect 23072 36332 23572 36360
rect 23072 36320 23078 36332
rect 23566 36320 23572 36332
rect 23624 36320 23630 36372
rect 23750 36320 23756 36372
rect 23808 36360 23814 36372
rect 24302 36360 24308 36372
rect 23808 36332 24308 36360
rect 23808 36320 23814 36332
rect 24302 36320 24308 36332
rect 24360 36320 24366 36372
rect 27893 36363 27951 36369
rect 27893 36329 27905 36363
rect 27939 36360 27951 36363
rect 28258 36360 28264 36372
rect 27939 36332 28264 36360
rect 27939 36329 27951 36332
rect 27893 36323 27951 36329
rect 28258 36320 28264 36332
rect 28316 36320 28322 36372
rect 29270 36320 29276 36372
rect 29328 36360 29334 36372
rect 30650 36360 30656 36372
rect 29328 36332 30656 36360
rect 29328 36320 29334 36332
rect 30650 36320 30656 36332
rect 30708 36320 30714 36372
rect 32214 36320 32220 36372
rect 32272 36320 32278 36372
rect 34054 36320 34060 36372
rect 34112 36320 34118 36372
rect 19978 36252 19984 36304
rect 20036 36292 20042 36304
rect 23934 36292 23940 36304
rect 20036 36264 23940 36292
rect 20036 36252 20042 36264
rect 23934 36252 23940 36264
rect 23992 36252 23998 36304
rect 24121 36295 24179 36301
rect 24121 36261 24133 36295
rect 24167 36292 24179 36295
rect 24486 36292 24492 36304
rect 24167 36264 24492 36292
rect 24167 36261 24179 36264
rect 24121 36255 24179 36261
rect 24486 36252 24492 36264
rect 24544 36252 24550 36304
rect 30006 36292 30012 36304
rect 25516 36264 30012 36292
rect 19334 36184 19340 36236
rect 19392 36224 19398 36236
rect 19797 36227 19855 36233
rect 19797 36224 19809 36227
rect 19392 36196 19809 36224
rect 19392 36184 19398 36196
rect 19797 36193 19809 36196
rect 19843 36193 19855 36227
rect 19797 36187 19855 36193
rect 22094 36184 22100 36236
rect 22152 36224 22158 36236
rect 23290 36224 23296 36236
rect 22152 36196 23296 36224
rect 22152 36184 22158 36196
rect 23290 36184 23296 36196
rect 23348 36224 23354 36236
rect 25516 36224 25544 36264
rect 30006 36252 30012 36264
rect 30064 36252 30070 36304
rect 32585 36295 32643 36301
rect 32585 36261 32597 36295
rect 32631 36261 32643 36295
rect 32585 36255 32643 36261
rect 27982 36224 27988 36236
rect 23348 36196 25544 36224
rect 23348 36184 23354 36196
rect 18509 36159 18567 36165
rect 18509 36156 18521 36159
rect 18104 36128 18521 36156
rect 18104 36116 18110 36128
rect 18509 36125 18521 36128
rect 18555 36125 18567 36159
rect 18509 36119 18567 36125
rect 18693 36159 18751 36165
rect 18693 36125 18705 36159
rect 18739 36125 18751 36159
rect 20170 36159 20228 36165
rect 20170 36156 20182 36159
rect 18693 36119 18751 36125
rect 18800 36128 20182 36156
rect 17328 36060 17540 36088
rect 17328 36020 17356 36060
rect 17586 36048 17592 36100
rect 17644 36088 17650 36100
rect 17681 36091 17739 36097
rect 17681 36088 17693 36091
rect 17644 36060 17693 36088
rect 17644 36048 17650 36060
rect 17681 36057 17693 36060
rect 17727 36057 17739 36091
rect 17880 36088 17908 36116
rect 18800 36088 18828 36128
rect 20170 36125 20182 36128
rect 20216 36125 20228 36159
rect 20170 36119 20228 36125
rect 22830 36116 22836 36168
rect 22888 36156 22894 36168
rect 23198 36156 23204 36168
rect 22888 36128 23204 36156
rect 22888 36116 22894 36128
rect 23198 36116 23204 36128
rect 23256 36156 23262 36168
rect 23569 36159 23627 36165
rect 23569 36156 23581 36159
rect 23256 36128 23581 36156
rect 23256 36116 23262 36128
rect 23569 36125 23581 36128
rect 23615 36125 23627 36159
rect 23569 36119 23627 36125
rect 23937 36159 23995 36165
rect 23937 36125 23949 36159
rect 23983 36156 23995 36159
rect 24578 36156 24584 36168
rect 23983 36128 24584 36156
rect 23983 36125 23995 36128
rect 23937 36119 23995 36125
rect 24578 36116 24584 36128
rect 24636 36116 24642 36168
rect 25516 36165 25544 36196
rect 27632 36196 27988 36224
rect 25501 36159 25559 36165
rect 25501 36125 25513 36159
rect 25547 36125 25559 36159
rect 25501 36119 25559 36125
rect 25777 36159 25835 36165
rect 25777 36125 25789 36159
rect 25823 36125 25835 36159
rect 25777 36119 25835 36125
rect 25869 36159 25927 36165
rect 25869 36125 25881 36159
rect 25915 36156 25927 36159
rect 25958 36156 25964 36168
rect 25915 36128 25964 36156
rect 25915 36125 25927 36128
rect 25869 36119 25927 36125
rect 17880 36060 18828 36088
rect 17681 36051 17739 36057
rect 19058 36048 19064 36100
rect 19116 36088 19122 36100
rect 19797 36091 19855 36097
rect 19797 36088 19809 36091
rect 19116 36060 19809 36088
rect 19116 36048 19122 36060
rect 19797 36057 19809 36060
rect 19843 36057 19855 36091
rect 19797 36051 19855 36057
rect 19978 36048 19984 36100
rect 20036 36048 20042 36100
rect 20073 36091 20131 36097
rect 20073 36057 20085 36091
rect 20119 36088 20131 36091
rect 20530 36088 20536 36100
rect 20119 36060 20536 36088
rect 20119 36057 20131 36060
rect 20073 36051 20131 36057
rect 20530 36048 20536 36060
rect 20588 36048 20594 36100
rect 21082 36048 21088 36100
rect 21140 36088 21146 36100
rect 23753 36091 23811 36097
rect 23753 36088 23765 36091
rect 21140 36060 23765 36088
rect 21140 36048 21146 36060
rect 23753 36057 23765 36060
rect 23799 36057 23811 36091
rect 23753 36051 23811 36057
rect 23845 36091 23903 36097
rect 23845 36057 23857 36091
rect 23891 36057 23903 36091
rect 23845 36051 23903 36057
rect 15948 35992 17356 36020
rect 17402 35980 17408 36032
rect 17460 35980 17466 36032
rect 18598 35980 18604 36032
rect 18656 35980 18662 36032
rect 22922 35980 22928 36032
rect 22980 36020 22986 36032
rect 23860 36020 23888 36051
rect 24946 36048 24952 36100
rect 25004 36088 25010 36100
rect 25685 36091 25743 36097
rect 25685 36088 25697 36091
rect 25004 36060 25697 36088
rect 25004 36048 25010 36060
rect 25685 36057 25697 36060
rect 25731 36057 25743 36091
rect 25685 36051 25743 36057
rect 25792 36088 25820 36119
rect 25958 36116 25964 36128
rect 26016 36116 26022 36168
rect 27246 36116 27252 36168
rect 27304 36116 27310 36168
rect 27338 36116 27344 36168
rect 27396 36156 27402 36168
rect 27632 36165 27660 36196
rect 27982 36184 27988 36196
rect 28040 36184 28046 36236
rect 28718 36184 28724 36236
rect 28776 36184 28782 36236
rect 27617 36159 27675 36165
rect 27396 36128 27441 36156
rect 27396 36116 27402 36128
rect 27617 36125 27629 36159
rect 27663 36125 27675 36159
rect 27617 36119 27675 36125
rect 27755 36159 27813 36165
rect 27755 36125 27767 36159
rect 27801 36156 27813 36159
rect 28258 36156 28264 36168
rect 27801 36128 28264 36156
rect 27801 36125 27813 36128
rect 27755 36119 27813 36125
rect 28258 36116 28264 36128
rect 28316 36116 28322 36168
rect 28534 36116 28540 36168
rect 28592 36116 28598 36168
rect 32033 36159 32091 36165
rect 32033 36125 32045 36159
rect 32079 36156 32091 36159
rect 32600 36156 32628 36255
rect 33137 36227 33195 36233
rect 33137 36224 33149 36227
rect 32079 36128 32628 36156
rect 32692 36196 33149 36224
rect 32079 36125 32091 36128
rect 32033 36119 32091 36125
rect 25792 36060 26188 36088
rect 25792 36020 25820 36060
rect 22980 35992 25820 36020
rect 22980 35980 22986 35992
rect 26050 35980 26056 36032
rect 26108 35980 26114 36032
rect 26160 36020 26188 36060
rect 26418 36048 26424 36100
rect 26476 36088 26482 36100
rect 27525 36091 27583 36097
rect 27525 36088 27537 36091
rect 26476 36060 27537 36088
rect 26476 36048 26482 36060
rect 27525 36057 27537 36060
rect 27571 36088 27583 36091
rect 29822 36088 29828 36100
rect 27571 36060 29828 36088
rect 27571 36057 27583 36060
rect 27525 36051 27583 36057
rect 29822 36048 29828 36060
rect 29880 36048 29886 36100
rect 30834 36048 30840 36100
rect 30892 36088 30898 36100
rect 32692 36088 32720 36196
rect 33137 36193 33149 36196
rect 33183 36193 33195 36227
rect 33137 36187 33195 36193
rect 33045 36159 33103 36165
rect 33045 36156 33057 36159
rect 30892 36060 32720 36088
rect 32784 36128 33057 36156
rect 30892 36048 30898 36060
rect 30742 36020 30748 36032
rect 26160 35992 30748 36020
rect 30742 35980 30748 35992
rect 30800 36020 30806 36032
rect 32784 36020 32812 36128
rect 33045 36125 33057 36128
rect 33091 36156 33103 36159
rect 34072 36156 34100 36320
rect 33091 36128 34100 36156
rect 33091 36125 33103 36128
rect 33045 36119 33103 36125
rect 30800 35992 32812 36020
rect 32953 36023 33011 36029
rect 30800 35980 30806 35992
rect 32953 35989 32965 36023
rect 32999 36020 33011 36023
rect 33134 36020 33140 36032
rect 32999 35992 33140 36020
rect 32999 35989 33011 35992
rect 32953 35983 33011 35989
rect 33134 35980 33140 35992
rect 33192 35980 33198 36032
rect 1104 35930 38272 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38272 35930
rect 1104 35856 38272 35878
rect 6270 35776 6276 35828
rect 6328 35816 6334 35828
rect 6549 35819 6607 35825
rect 6549 35816 6561 35819
rect 6328 35788 6561 35816
rect 6328 35776 6334 35788
rect 6549 35785 6561 35788
rect 6595 35785 6607 35819
rect 6549 35779 6607 35785
rect 7653 35819 7711 35825
rect 7653 35785 7665 35819
rect 7699 35816 7711 35819
rect 7742 35816 7748 35828
rect 7699 35788 7748 35816
rect 7699 35785 7711 35788
rect 7653 35779 7711 35785
rect 7742 35776 7748 35788
rect 7800 35816 7806 35828
rect 8110 35816 8116 35828
rect 7800 35788 8116 35816
rect 7800 35776 7806 35788
rect 8110 35776 8116 35788
rect 8168 35776 8174 35828
rect 9122 35776 9128 35828
rect 9180 35816 9186 35828
rect 12894 35816 12900 35828
rect 9180 35788 12900 35816
rect 9180 35776 9186 35788
rect 12894 35776 12900 35788
rect 12952 35776 12958 35828
rect 13354 35816 13360 35828
rect 13188 35788 13360 35816
rect 9493 35751 9551 35757
rect 9493 35717 9505 35751
rect 9539 35748 9551 35751
rect 9582 35748 9588 35760
rect 9539 35720 9588 35748
rect 9539 35717 9551 35720
rect 9493 35711 9551 35717
rect 9582 35708 9588 35720
rect 9640 35708 9646 35760
rect 10226 35708 10232 35760
rect 10284 35708 10290 35760
rect 11146 35708 11152 35760
rect 11204 35748 11210 35760
rect 12986 35748 12992 35760
rect 11204 35720 12992 35748
rect 11204 35708 11210 35720
rect 12986 35708 12992 35720
rect 13044 35708 13050 35760
rect 6733 35683 6791 35689
rect 6733 35649 6745 35683
rect 6779 35680 6791 35683
rect 7745 35683 7803 35689
rect 6779 35652 6914 35680
rect 6779 35649 6791 35652
rect 6733 35643 6791 35649
rect 6886 35544 6914 35652
rect 7745 35649 7757 35683
rect 7791 35680 7803 35683
rect 9125 35683 9183 35689
rect 7791 35652 8248 35680
rect 7791 35649 7803 35652
rect 7745 35643 7803 35649
rect 8220 35624 8248 35652
rect 9125 35649 9137 35683
rect 9171 35649 9183 35683
rect 9125 35643 9183 35649
rect 7466 35572 7472 35624
rect 7524 35612 7530 35624
rect 7837 35615 7895 35621
rect 7837 35612 7849 35615
rect 7524 35584 7849 35612
rect 7524 35572 7530 35584
rect 7837 35581 7849 35584
rect 7883 35581 7895 35615
rect 7837 35575 7895 35581
rect 8202 35572 8208 35624
rect 8260 35572 8266 35624
rect 8294 35572 8300 35624
rect 8352 35572 8358 35624
rect 9140 35612 9168 35643
rect 9214 35640 9220 35692
rect 9272 35640 9278 35692
rect 13081 35683 13139 35689
rect 13081 35649 13093 35683
rect 13127 35680 13139 35683
rect 13188 35680 13216 35788
rect 13354 35776 13360 35788
rect 13412 35816 13418 35828
rect 13633 35819 13691 35825
rect 13633 35816 13645 35819
rect 13412 35788 13645 35816
rect 13412 35776 13418 35788
rect 13633 35785 13645 35788
rect 13679 35785 13691 35819
rect 13633 35779 13691 35785
rect 13909 35819 13967 35825
rect 13909 35785 13921 35819
rect 13955 35816 13967 35819
rect 14274 35816 14280 35828
rect 13955 35788 14280 35816
rect 13955 35785 13967 35788
rect 13909 35779 13967 35785
rect 14274 35776 14280 35788
rect 14332 35776 14338 35828
rect 23290 35816 23296 35828
rect 23124 35788 23296 35816
rect 13265 35751 13323 35757
rect 13265 35717 13277 35751
rect 13311 35748 13323 35751
rect 14001 35751 14059 35757
rect 14001 35748 14013 35751
rect 13311 35720 14013 35748
rect 13311 35717 13323 35720
rect 13265 35711 13323 35717
rect 14001 35717 14013 35720
rect 14047 35717 14059 35751
rect 14001 35711 14059 35717
rect 18598 35708 18604 35760
rect 18656 35748 18662 35760
rect 19061 35751 19119 35757
rect 19061 35748 19073 35751
rect 18656 35720 19073 35748
rect 18656 35708 18662 35720
rect 19061 35717 19073 35720
rect 19107 35717 19119 35751
rect 19061 35711 19119 35717
rect 20438 35708 20444 35760
rect 20496 35748 20502 35760
rect 21085 35751 21143 35757
rect 21085 35748 21097 35751
rect 20496 35720 21097 35748
rect 20496 35708 20502 35720
rect 21085 35717 21097 35720
rect 21131 35717 21143 35751
rect 21085 35711 21143 35717
rect 22186 35708 22192 35760
rect 22244 35708 22250 35760
rect 13127 35652 13216 35680
rect 13127 35649 13139 35652
rect 13081 35643 13139 35649
rect 13538 35640 13544 35692
rect 13596 35640 13602 35692
rect 13722 35640 13728 35692
rect 13780 35640 13786 35692
rect 14829 35683 14887 35689
rect 14829 35649 14841 35683
rect 14875 35680 14887 35683
rect 14875 35652 18000 35680
rect 14875 35649 14887 35652
rect 14829 35643 14887 35649
rect 9490 35612 9496 35624
rect 9140 35584 9496 35612
rect 9490 35572 9496 35584
rect 9548 35572 9554 35624
rect 12897 35615 12955 35621
rect 12897 35581 12909 35615
rect 12943 35612 12955 35615
rect 13556 35612 13584 35640
rect 12943 35584 13584 35612
rect 12943 35581 12955 35584
rect 12897 35575 12955 35581
rect 13630 35572 13636 35624
rect 13688 35612 13694 35624
rect 14844 35612 14872 35643
rect 17972 35624 18000 35652
rect 18874 35640 18880 35692
rect 18932 35640 18938 35692
rect 18969 35683 19027 35689
rect 18969 35649 18981 35683
rect 19015 35649 19027 35683
rect 18969 35643 19027 35649
rect 19199 35683 19257 35689
rect 19199 35649 19211 35683
rect 19245 35680 19257 35683
rect 19978 35680 19984 35692
rect 19245 35652 19984 35680
rect 19245 35649 19257 35652
rect 19199 35643 19257 35649
rect 13688 35584 14872 35612
rect 13688 35572 13694 35584
rect 16206 35572 16212 35624
rect 16264 35572 16270 35624
rect 17954 35572 17960 35624
rect 18012 35572 18018 35624
rect 7285 35547 7343 35553
rect 7285 35544 7297 35547
rect 6886 35516 7297 35544
rect 7285 35513 7297 35516
rect 7331 35513 7343 35547
rect 7285 35507 7343 35513
rect 11330 35504 11336 35556
rect 11388 35544 11394 35556
rect 13357 35547 13415 35553
rect 13357 35544 13369 35547
rect 11388 35516 13369 35544
rect 11388 35504 11394 35516
rect 13357 35513 13369 35516
rect 13403 35544 13415 35547
rect 16224 35544 16252 35572
rect 13403 35516 16252 35544
rect 18984 35544 19012 35643
rect 19978 35640 19984 35652
rect 20036 35640 20042 35692
rect 20070 35640 20076 35692
rect 20128 35680 20134 35692
rect 20993 35683 21051 35689
rect 20993 35680 21005 35683
rect 20128 35652 21005 35680
rect 20128 35640 20134 35652
rect 20993 35649 21005 35652
rect 21039 35649 21051 35683
rect 20993 35643 21051 35649
rect 21174 35640 21180 35692
rect 21232 35640 21238 35692
rect 22094 35689 22100 35692
rect 21361 35683 21419 35689
rect 21361 35649 21373 35683
rect 21407 35680 21419 35683
rect 21913 35683 21971 35689
rect 21913 35680 21925 35683
rect 21407 35652 21925 35680
rect 21407 35649 21419 35652
rect 21361 35643 21419 35649
rect 21913 35649 21925 35652
rect 21959 35649 21971 35683
rect 21913 35643 21971 35649
rect 22061 35683 22100 35689
rect 22061 35649 22073 35683
rect 22061 35643 22100 35649
rect 22094 35640 22100 35643
rect 22152 35640 22158 35692
rect 22278 35680 22284 35692
rect 22239 35652 22284 35680
rect 22278 35640 22284 35652
rect 22336 35640 22342 35692
rect 22370 35640 22376 35692
rect 22428 35689 22434 35692
rect 22428 35680 22436 35689
rect 22428 35652 22473 35680
rect 22428 35643 22436 35652
rect 22428 35640 22434 35643
rect 22554 35640 22560 35692
rect 22612 35640 22618 35692
rect 22830 35640 22836 35692
rect 22888 35640 22894 35692
rect 22922 35640 22928 35692
rect 22980 35680 22986 35692
rect 23124 35689 23152 35788
rect 23290 35776 23296 35788
rect 23348 35776 23354 35828
rect 23658 35776 23664 35828
rect 23716 35816 23722 35828
rect 25958 35816 25964 35828
rect 23716 35788 24164 35816
rect 23716 35776 23722 35788
rect 23198 35708 23204 35760
rect 23256 35708 23262 35760
rect 23845 35751 23903 35757
rect 23845 35717 23857 35751
rect 23891 35748 23903 35751
rect 24026 35748 24032 35760
rect 23891 35720 24032 35748
rect 23891 35717 23903 35720
rect 23845 35711 23903 35717
rect 24026 35708 24032 35720
rect 24084 35708 24090 35760
rect 23109 35683 23167 35689
rect 22980 35652 23025 35680
rect 22980 35640 22986 35652
rect 23109 35649 23121 35683
rect 23155 35649 23167 35683
rect 23298 35683 23356 35689
rect 23298 35680 23310 35683
rect 23109 35643 23167 35649
rect 23216 35652 23310 35680
rect 19337 35615 19395 35621
rect 19337 35581 19349 35615
rect 19383 35612 19395 35615
rect 21450 35612 21456 35624
rect 19383 35584 21456 35612
rect 19383 35581 19395 35584
rect 19337 35575 19395 35581
rect 21450 35572 21456 35584
rect 21508 35572 21514 35624
rect 22572 35612 22600 35640
rect 22738 35612 22744 35624
rect 22572 35584 22744 35612
rect 22738 35572 22744 35584
rect 22796 35612 22802 35624
rect 23216 35612 23244 35652
rect 23298 35649 23310 35652
rect 23344 35649 23356 35683
rect 23298 35643 23356 35649
rect 23750 35640 23756 35692
rect 23808 35640 23814 35692
rect 24136 35689 24164 35788
rect 25240 35788 25964 35816
rect 25130 35708 25136 35760
rect 25188 35708 25194 35760
rect 23937 35683 23995 35689
rect 23937 35649 23949 35683
rect 23983 35649 23995 35683
rect 23937 35643 23995 35649
rect 24121 35683 24179 35689
rect 24121 35649 24133 35683
rect 24167 35649 24179 35683
rect 24121 35643 24179 35649
rect 22796 35584 23244 35612
rect 22796 35572 22802 35584
rect 23842 35572 23848 35624
rect 23900 35612 23906 35624
rect 23952 35612 23980 35643
rect 23900 35584 23980 35612
rect 24136 35612 24164 35643
rect 24854 35640 24860 35692
rect 24912 35640 24918 35692
rect 24946 35640 24952 35692
rect 25004 35680 25010 35692
rect 25240 35689 25268 35788
rect 25958 35776 25964 35788
rect 26016 35776 26022 35828
rect 26050 35776 26056 35828
rect 26108 35776 26114 35828
rect 27798 35776 27804 35828
rect 27856 35816 27862 35828
rect 29181 35819 29239 35825
rect 29181 35816 29193 35819
rect 27856 35788 29193 35816
rect 27856 35776 27862 35788
rect 29181 35785 29193 35788
rect 29227 35785 29239 35819
rect 29181 35779 29239 35785
rect 29564 35788 30696 35816
rect 26068 35748 26096 35776
rect 25332 35720 25820 35748
rect 25041 35683 25099 35689
rect 25041 35680 25053 35683
rect 25004 35652 25053 35680
rect 25004 35640 25010 35652
rect 25041 35649 25053 35652
rect 25087 35649 25099 35683
rect 25041 35643 25099 35649
rect 25225 35683 25283 35689
rect 25225 35649 25237 35683
rect 25271 35649 25283 35683
rect 25225 35643 25283 35649
rect 25332 35612 25360 35720
rect 25406 35640 25412 35692
rect 25464 35680 25470 35692
rect 25792 35689 25820 35720
rect 25976 35720 26096 35748
rect 25685 35683 25743 35689
rect 25685 35680 25697 35683
rect 25464 35652 25697 35680
rect 25464 35640 25470 35652
rect 25685 35649 25697 35652
rect 25731 35649 25743 35683
rect 25685 35643 25743 35649
rect 25777 35683 25835 35689
rect 25777 35649 25789 35683
rect 25823 35680 25835 35683
rect 25866 35680 25872 35692
rect 25823 35652 25872 35680
rect 25823 35649 25835 35652
rect 25777 35643 25835 35649
rect 25866 35640 25872 35652
rect 25924 35640 25930 35692
rect 25976 35689 26004 35720
rect 28718 35708 28724 35760
rect 28776 35708 28782 35760
rect 25961 35683 26019 35689
rect 25961 35649 25973 35683
rect 26007 35649 26019 35683
rect 25961 35643 26019 35649
rect 26050 35640 26056 35692
rect 26108 35680 26114 35692
rect 26145 35683 26203 35689
rect 26145 35680 26157 35683
rect 26108 35652 26157 35680
rect 26108 35640 26114 35652
rect 26145 35649 26157 35652
rect 26191 35649 26203 35683
rect 26145 35643 26203 35649
rect 26237 35683 26295 35689
rect 26237 35649 26249 35683
rect 26283 35649 26295 35683
rect 26237 35643 26295 35649
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35649 26479 35683
rect 26421 35643 26479 35649
rect 26252 35612 26280 35643
rect 24136 35584 25360 35612
rect 25792 35584 26280 35612
rect 26436 35612 26464 35643
rect 26510 35640 26516 35692
rect 26568 35640 26574 35692
rect 27338 35640 27344 35692
rect 27396 35640 27402 35692
rect 29564 35680 29592 35788
rect 30466 35748 30472 35760
rect 29656 35720 30472 35748
rect 29656 35689 29684 35720
rect 30466 35708 30472 35720
rect 30524 35708 30530 35760
rect 28966 35652 29592 35680
rect 29641 35683 29699 35689
rect 27356 35612 27384 35640
rect 26436 35584 27384 35612
rect 23900 35572 23906 35584
rect 20809 35547 20867 35553
rect 18984 35516 19380 35544
rect 13403 35513 13415 35516
rect 13357 35507 13415 35513
rect 19352 35488 19380 35516
rect 20809 35513 20821 35547
rect 20855 35544 20867 35547
rect 20990 35544 20996 35556
rect 20855 35516 20996 35544
rect 20855 35513 20867 35516
rect 20809 35507 20867 35513
rect 20990 35504 20996 35516
rect 21048 35504 21054 35556
rect 22557 35547 22615 35553
rect 22557 35513 22569 35547
rect 22603 35544 22615 35547
rect 23658 35544 23664 35556
rect 22603 35516 23664 35544
rect 22603 35513 22615 35516
rect 22557 35507 22615 35513
rect 23658 35504 23664 35516
rect 23716 35504 23722 35556
rect 25409 35547 25467 35553
rect 25409 35513 25421 35547
rect 25455 35544 25467 35547
rect 25792 35544 25820 35584
rect 27430 35572 27436 35624
rect 27488 35572 27494 35624
rect 27709 35615 27767 35621
rect 27709 35581 27721 35615
rect 27755 35612 27767 35615
rect 28166 35612 28172 35624
rect 27755 35584 28172 35612
rect 27755 35581 27767 35584
rect 27709 35575 27767 35581
rect 28166 35572 28172 35584
rect 28224 35572 28230 35624
rect 28258 35572 28264 35624
rect 28316 35612 28322 35624
rect 28442 35612 28448 35624
rect 28316 35584 28448 35612
rect 28316 35572 28322 35584
rect 28442 35572 28448 35584
rect 28500 35612 28506 35624
rect 28966 35612 28994 35652
rect 29641 35649 29653 35683
rect 29687 35649 29699 35683
rect 29641 35643 29699 35649
rect 29734 35683 29792 35689
rect 29734 35649 29746 35683
rect 29780 35649 29792 35683
rect 29734 35643 29792 35649
rect 29748 35612 29776 35643
rect 29822 35640 29828 35692
rect 29880 35680 29886 35692
rect 29917 35683 29975 35689
rect 29917 35680 29929 35683
rect 29880 35652 29929 35680
rect 29880 35640 29886 35652
rect 29917 35649 29929 35652
rect 29963 35649 29975 35683
rect 29917 35643 29975 35649
rect 30006 35640 30012 35692
rect 30064 35640 30070 35692
rect 30106 35683 30164 35689
rect 30106 35649 30118 35683
rect 30152 35649 30164 35683
rect 30561 35683 30619 35689
rect 30561 35680 30573 35683
rect 30106 35643 30164 35649
rect 30300 35652 30573 35680
rect 30116 35612 30144 35643
rect 28500 35584 28994 35612
rect 29656 35584 29776 35612
rect 29932 35584 30144 35612
rect 28500 35572 28506 35584
rect 25455 35516 25820 35544
rect 25455 35513 25467 35516
rect 25409 35507 25467 35513
rect 25866 35504 25872 35556
rect 25924 35544 25930 35556
rect 25924 35516 27568 35544
rect 25924 35504 25930 35516
rect 10962 35436 10968 35488
rect 11020 35476 11026 35488
rect 12526 35476 12532 35488
rect 11020 35448 12532 35476
rect 11020 35436 11026 35448
rect 12526 35436 12532 35448
rect 12584 35436 12590 35488
rect 18690 35436 18696 35488
rect 18748 35436 18754 35488
rect 19334 35436 19340 35488
rect 19392 35436 19398 35488
rect 23474 35436 23480 35488
rect 23532 35436 23538 35488
rect 23569 35479 23627 35485
rect 23569 35445 23581 35479
rect 23615 35476 23627 35479
rect 23934 35476 23940 35488
rect 23615 35448 23940 35476
rect 23615 35445 23627 35448
rect 23569 35439 23627 35445
rect 23934 35436 23940 35448
rect 23992 35436 23998 35488
rect 25498 35436 25504 35488
rect 25556 35436 25562 35488
rect 26602 35436 26608 35488
rect 26660 35476 26666 35488
rect 26697 35479 26755 35485
rect 26697 35476 26709 35479
rect 26660 35448 26709 35476
rect 26660 35436 26666 35448
rect 26697 35445 26709 35448
rect 26743 35445 26755 35479
rect 27540 35476 27568 35516
rect 29656 35488 29684 35584
rect 29932 35488 29960 35584
rect 30300 35553 30328 35652
rect 30561 35649 30573 35652
rect 30607 35649 30619 35683
rect 30668 35680 30696 35788
rect 30742 35776 30748 35828
rect 30800 35776 30806 35828
rect 32582 35708 32588 35760
rect 32640 35708 32646 35760
rect 30837 35683 30895 35689
rect 30837 35680 30849 35683
rect 30668 35652 30849 35680
rect 30561 35643 30619 35649
rect 30837 35649 30849 35652
rect 30883 35649 30895 35683
rect 30837 35643 30895 35649
rect 30852 35612 30880 35643
rect 31386 35640 31392 35692
rect 31444 35640 31450 35692
rect 32600 35680 32628 35708
rect 32953 35683 33011 35689
rect 32953 35680 32965 35683
rect 32600 35652 32965 35680
rect 32953 35649 32965 35652
rect 32999 35649 33011 35683
rect 32953 35643 33011 35649
rect 33502 35640 33508 35692
rect 33560 35640 33566 35692
rect 31478 35612 31484 35624
rect 30852 35584 31484 35612
rect 31478 35572 31484 35584
rect 31536 35572 31542 35624
rect 30285 35547 30343 35553
rect 30285 35513 30297 35547
rect 30331 35513 30343 35547
rect 30285 35507 30343 35513
rect 29638 35476 29644 35488
rect 27540 35448 29644 35476
rect 26697 35439 26755 35445
rect 29638 35436 29644 35448
rect 29696 35436 29702 35488
rect 29914 35436 29920 35488
rect 29972 35436 29978 35488
rect 30098 35436 30104 35488
rect 30156 35476 30162 35488
rect 30377 35479 30435 35485
rect 30377 35476 30389 35479
rect 30156 35448 30389 35476
rect 30156 35436 30162 35448
rect 30377 35445 30389 35448
rect 30423 35445 30435 35479
rect 30377 35439 30435 35445
rect 31018 35436 31024 35488
rect 31076 35476 31082 35488
rect 31205 35479 31263 35485
rect 31205 35476 31217 35479
rect 31076 35448 31217 35476
rect 31076 35436 31082 35448
rect 31205 35445 31217 35448
rect 31251 35445 31263 35479
rect 31205 35439 31263 35445
rect 32766 35436 32772 35488
rect 32824 35476 32830 35488
rect 32861 35479 32919 35485
rect 32861 35476 32873 35479
rect 32824 35448 32873 35476
rect 32824 35436 32830 35448
rect 32861 35445 32873 35448
rect 32907 35445 32919 35479
rect 32861 35439 32919 35445
rect 33318 35436 33324 35488
rect 33376 35436 33382 35488
rect 1104 35386 38272 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38272 35386
rect 1104 35312 38272 35334
rect 9493 35275 9551 35281
rect 9493 35241 9505 35275
rect 9539 35272 9551 35275
rect 9766 35272 9772 35284
rect 9539 35244 9772 35272
rect 9539 35241 9551 35244
rect 9493 35235 9551 35241
rect 9766 35232 9772 35244
rect 9824 35232 9830 35284
rect 10962 35232 10968 35284
rect 11020 35232 11026 35284
rect 17497 35275 17555 35281
rect 17497 35241 17509 35275
rect 17543 35272 17555 35275
rect 18874 35272 18880 35284
rect 17543 35244 18880 35272
rect 17543 35241 17555 35244
rect 17497 35235 17555 35241
rect 18874 35232 18880 35244
rect 18932 35232 18938 35284
rect 23474 35232 23480 35284
rect 23532 35232 23538 35284
rect 23934 35232 23940 35284
rect 23992 35232 23998 35284
rect 25406 35232 25412 35284
rect 25464 35272 25470 35284
rect 26510 35272 26516 35284
rect 25464 35244 26516 35272
rect 25464 35232 25470 35244
rect 26510 35232 26516 35244
rect 26568 35232 26574 35284
rect 28166 35232 28172 35284
rect 28224 35232 28230 35284
rect 28350 35232 28356 35284
rect 28408 35272 28414 35284
rect 29914 35272 29920 35284
rect 28408 35244 29920 35272
rect 28408 35232 28414 35244
rect 29914 35232 29920 35244
rect 29972 35232 29978 35284
rect 32766 35232 32772 35284
rect 32824 35232 32830 35284
rect 9858 35164 9864 35216
rect 9916 35204 9922 35216
rect 10778 35204 10784 35216
rect 9916 35176 10784 35204
rect 9916 35164 9922 35176
rect 7190 35136 7196 35148
rect 6656 35108 7196 35136
rect 6656 35077 6684 35108
rect 7190 35096 7196 35108
rect 7248 35096 7254 35148
rect 10060 35145 10088 35176
rect 10778 35164 10784 35176
rect 10836 35164 10842 35216
rect 9953 35139 10011 35145
rect 9953 35136 9965 35139
rect 8220 35108 9965 35136
rect 8220 35080 8248 35108
rect 9953 35105 9965 35108
rect 9999 35105 10011 35139
rect 9953 35099 10011 35105
rect 10045 35139 10103 35145
rect 10045 35105 10057 35139
rect 10091 35105 10103 35139
rect 10045 35099 10103 35105
rect 6641 35071 6699 35077
rect 6641 35037 6653 35071
rect 6687 35037 6699 35071
rect 6641 35031 6699 35037
rect 6733 35071 6791 35077
rect 6733 35037 6745 35071
rect 6779 35068 6791 35071
rect 6917 35071 6975 35077
rect 6917 35068 6929 35071
rect 6779 35040 6929 35068
rect 6779 35037 6791 35040
rect 6733 35031 6791 35037
rect 6917 35037 6929 35040
rect 6963 35037 6975 35071
rect 6917 35031 6975 35037
rect 8202 35028 8208 35080
rect 8260 35028 8266 35080
rect 8294 35028 8300 35080
rect 8352 35028 8358 35080
rect 9861 35071 9919 35077
rect 9861 35037 9873 35071
rect 9907 35068 9919 35071
rect 10980 35068 11008 35232
rect 15102 35096 15108 35148
rect 15160 35136 15166 35148
rect 18782 35136 18788 35148
rect 15160 35108 18788 35136
rect 15160 35096 15166 35108
rect 18782 35096 18788 35108
rect 18840 35096 18846 35148
rect 20990 35096 20996 35148
rect 21048 35136 21054 35148
rect 22554 35136 22560 35148
rect 21048 35108 22560 35136
rect 21048 35096 21054 35108
rect 22554 35096 22560 35108
rect 22612 35096 22618 35148
rect 23492 35136 23520 35232
rect 23952 35204 23980 35232
rect 23860 35176 23980 35204
rect 23569 35139 23627 35145
rect 23569 35136 23581 35139
rect 23492 35108 23581 35136
rect 23569 35105 23581 35108
rect 23615 35105 23627 35139
rect 23569 35099 23627 35105
rect 23658 35096 23664 35148
rect 23716 35096 23722 35148
rect 9907 35040 11008 35068
rect 9907 35037 9919 35040
rect 9861 35031 9919 35037
rect 17310 35028 17316 35080
rect 17368 35028 17374 35080
rect 20806 35028 20812 35080
rect 20864 35068 20870 35080
rect 23293 35071 23351 35077
rect 23293 35068 23305 35071
rect 20864 35040 23305 35068
rect 20864 35028 20870 35040
rect 23293 35037 23305 35040
rect 23339 35037 23351 35071
rect 23293 35031 23351 35037
rect 23477 35071 23535 35077
rect 23477 35037 23489 35071
rect 23523 35068 23535 35071
rect 23753 35071 23811 35077
rect 23523 35040 23704 35068
rect 23523 35037 23535 35040
rect 23477 35031 23535 35037
rect 7190 34960 7196 35012
rect 7248 34960 7254 35012
rect 16114 34960 16120 35012
rect 16172 35000 16178 35012
rect 18138 35000 18144 35012
rect 16172 34972 18144 35000
rect 16172 34960 16178 34972
rect 18138 34960 18144 34972
rect 18196 34960 18202 35012
rect 23566 35000 23572 35012
rect 22296 34972 23572 35000
rect 22296 34944 22324 34972
rect 23566 34960 23572 34972
rect 23624 34960 23630 35012
rect 23676 35000 23704 35040
rect 23753 35037 23765 35071
rect 23799 35068 23811 35071
rect 23860 35068 23888 35176
rect 24854 35164 24860 35216
rect 24912 35204 24918 35216
rect 26142 35204 26148 35216
rect 24912 35176 26148 35204
rect 24912 35164 24918 35176
rect 26068 35145 26096 35176
rect 26142 35164 26148 35176
rect 26200 35164 26206 35216
rect 26252 35176 27384 35204
rect 26053 35139 26111 35145
rect 23799 35040 23888 35068
rect 23952 35108 25728 35136
rect 23799 35037 23811 35040
rect 23753 35031 23811 35037
rect 23952 35000 23980 35108
rect 25314 35028 25320 35080
rect 25372 35028 25378 35080
rect 25498 35028 25504 35080
rect 25556 35028 25562 35080
rect 25700 35077 25728 35108
rect 26053 35105 26065 35139
rect 26099 35105 26111 35139
rect 26053 35099 26111 35105
rect 25593 35071 25651 35077
rect 25593 35037 25605 35071
rect 25639 35037 25651 35071
rect 25593 35031 25651 35037
rect 25685 35071 25743 35077
rect 25685 35037 25697 35071
rect 25731 35068 25743 35071
rect 26252 35068 26280 35176
rect 26602 35136 26608 35148
rect 26528 35108 26608 35136
rect 25731 35040 26280 35068
rect 25731 35037 25743 35040
rect 25685 35031 25743 35037
rect 23676 34972 23980 35000
rect 25608 35000 25636 35031
rect 26326 35028 26332 35080
rect 26384 35028 26390 35080
rect 26528 35077 26556 35108
rect 26602 35096 26608 35108
rect 26660 35096 26666 35148
rect 27356 35080 27384 35176
rect 28074 35164 28080 35216
rect 28132 35164 28138 35216
rect 29546 35164 29552 35216
rect 29604 35164 29610 35216
rect 27525 35139 27583 35145
rect 27525 35105 27537 35139
rect 27571 35136 27583 35139
rect 27571 35108 27844 35136
rect 27571 35105 27583 35108
rect 27525 35099 27583 35105
rect 26421 35071 26479 35077
rect 26421 35037 26433 35071
rect 26467 35037 26479 35071
rect 26421 35031 26479 35037
rect 26513 35071 26571 35077
rect 26513 35037 26525 35071
rect 26559 35037 26571 35071
rect 26513 35031 26571 35037
rect 26436 35000 26464 35031
rect 26694 35028 26700 35080
rect 26752 35028 26758 35080
rect 27338 35028 27344 35080
rect 27396 35028 27402 35080
rect 27614 35028 27620 35080
rect 27672 35068 27678 35080
rect 27709 35071 27767 35077
rect 27709 35068 27721 35071
rect 27672 35040 27721 35068
rect 27672 35028 27678 35040
rect 27709 35037 27721 35040
rect 27755 35037 27767 35071
rect 27709 35031 27767 35037
rect 26786 35000 26792 35012
rect 25608 34972 26792 35000
rect 26786 34960 26792 34972
rect 26844 34960 26850 35012
rect 27816 35000 27844 35108
rect 27908 35108 28948 35136
rect 27908 35080 27936 35108
rect 27890 35028 27896 35080
rect 27948 35028 27954 35080
rect 28074 35028 28080 35080
rect 28132 35068 28138 35080
rect 28920 35077 28948 35108
rect 28353 35071 28411 35077
rect 28353 35068 28365 35071
rect 28132 35040 28365 35068
rect 28132 35028 28138 35040
rect 28353 35037 28365 35040
rect 28399 35037 28411 35071
rect 28905 35071 28963 35077
rect 28905 35068 28917 35071
rect 28863 35040 28917 35068
rect 28353 35031 28411 35037
rect 28905 35037 28917 35040
rect 28951 35068 28963 35071
rect 29564 35068 29592 35164
rect 30929 35139 30987 35145
rect 30929 35105 30941 35139
rect 30975 35136 30987 35139
rect 31018 35136 31024 35148
rect 30975 35108 31024 35136
rect 30975 35105 30987 35108
rect 30929 35099 30987 35105
rect 31018 35096 31024 35108
rect 31076 35096 31082 35148
rect 32677 35139 32735 35145
rect 32677 35105 32689 35139
rect 32723 35136 32735 35139
rect 32784 35136 32812 35232
rect 32723 35108 32812 35136
rect 32953 35139 33011 35145
rect 32723 35105 32735 35108
rect 32677 35099 32735 35105
rect 32953 35105 32965 35139
rect 32999 35136 33011 35139
rect 33318 35136 33324 35148
rect 32999 35108 33324 35136
rect 32999 35105 33011 35108
rect 32953 35099 33011 35105
rect 33318 35096 33324 35108
rect 33376 35096 33382 35148
rect 33410 35096 33416 35148
rect 33468 35136 33474 35148
rect 33686 35136 33692 35148
rect 33468 35108 33692 35136
rect 33468 35096 33474 35108
rect 33686 35096 33692 35108
rect 33744 35096 33750 35148
rect 28951 35040 29592 35068
rect 28951 35037 28963 35040
rect 28905 35031 28963 35037
rect 30374 35028 30380 35080
rect 30432 35028 30438 35080
rect 30469 35071 30527 35077
rect 30469 35037 30481 35071
rect 30515 35068 30527 35071
rect 30653 35071 30711 35077
rect 30653 35068 30665 35071
rect 30515 35040 30665 35068
rect 30515 35037 30527 35040
rect 30469 35031 30527 35037
rect 30653 35037 30665 35040
rect 30699 35037 30711 35071
rect 30653 35031 30711 35037
rect 30834 35000 30840 35012
rect 27816 34972 30840 35000
rect 30834 34960 30840 34972
rect 30892 34960 30898 35012
rect 32490 35000 32496 35012
rect 32154 34972 32496 35000
rect 32490 34960 32496 34972
rect 32548 35000 32554 35012
rect 33410 35000 33416 35012
rect 32548 34972 33416 35000
rect 32548 34960 32554 34972
rect 33410 34960 33416 34972
rect 33468 34960 33474 35012
rect 8662 34892 8668 34944
rect 8720 34892 8726 34944
rect 13078 34892 13084 34944
rect 13136 34932 13142 34944
rect 20714 34932 20720 34944
rect 13136 34904 20720 34932
rect 13136 34892 13142 34904
rect 20714 34892 20720 34904
rect 20772 34892 20778 34944
rect 22278 34892 22284 34944
rect 22336 34892 22342 34944
rect 22922 34892 22928 34944
rect 22980 34932 22986 34944
rect 23842 34932 23848 34944
rect 22980 34904 23848 34932
rect 22980 34892 22986 34904
rect 23842 34892 23848 34904
rect 23900 34892 23906 34944
rect 23934 34892 23940 34944
rect 23992 34892 23998 34944
rect 25222 34892 25228 34944
rect 25280 34932 25286 34944
rect 25590 34932 25596 34944
rect 25280 34904 25596 34932
rect 25280 34892 25286 34904
rect 25590 34892 25596 34904
rect 25648 34932 25654 34944
rect 25961 34935 26019 34941
rect 25961 34932 25973 34935
rect 25648 34904 25973 34932
rect 25648 34892 25654 34904
rect 25961 34901 25973 34904
rect 26007 34901 26019 34935
rect 25961 34895 26019 34901
rect 27617 34935 27675 34941
rect 27617 34901 27629 34935
rect 27663 34932 27675 34935
rect 27798 34932 27804 34944
rect 27663 34904 27804 34932
rect 27663 34901 27675 34904
rect 27617 34895 27675 34901
rect 27798 34892 27804 34904
rect 27856 34892 27862 34944
rect 28810 34892 28816 34944
rect 28868 34892 28874 34944
rect 31662 34892 31668 34944
rect 31720 34932 31726 34944
rect 32401 34935 32459 34941
rect 32401 34932 32413 34935
rect 31720 34904 32413 34932
rect 31720 34892 31726 34904
rect 32401 34901 32413 34904
rect 32447 34901 32459 34935
rect 32401 34895 32459 34901
rect 33318 34892 33324 34944
rect 33376 34932 33382 34944
rect 34425 34935 34483 34941
rect 34425 34932 34437 34935
rect 33376 34904 34437 34932
rect 33376 34892 33382 34904
rect 34425 34901 34437 34904
rect 34471 34901 34483 34935
rect 34425 34895 34483 34901
rect 1104 34842 38272 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38272 34842
rect 1104 34768 38272 34790
rect 7190 34688 7196 34740
rect 7248 34728 7254 34740
rect 7653 34731 7711 34737
rect 7653 34728 7665 34731
rect 7248 34700 7665 34728
rect 7248 34688 7254 34700
rect 7653 34697 7665 34700
rect 7699 34697 7711 34731
rect 7653 34691 7711 34697
rect 7929 34731 7987 34737
rect 7929 34697 7941 34731
rect 7975 34697 7987 34731
rect 7929 34691 7987 34697
rect 5534 34552 5540 34604
rect 5592 34592 5598 34604
rect 5629 34595 5687 34601
rect 5629 34592 5641 34595
rect 5592 34564 5641 34592
rect 5592 34552 5598 34564
rect 5629 34561 5641 34564
rect 5675 34561 5687 34595
rect 5629 34555 5687 34561
rect 7837 34595 7895 34601
rect 7837 34561 7849 34595
rect 7883 34592 7895 34595
rect 7944 34592 7972 34691
rect 11698 34688 11704 34740
rect 11756 34728 11762 34740
rect 13630 34728 13636 34740
rect 11756 34700 13636 34728
rect 11756 34688 11762 34700
rect 13630 34688 13636 34700
rect 13688 34688 13694 34740
rect 16853 34731 16911 34737
rect 16853 34697 16865 34731
rect 16899 34728 16911 34731
rect 17310 34728 17316 34740
rect 16899 34700 17316 34728
rect 16899 34697 16911 34700
rect 16853 34691 16911 34697
rect 17310 34688 17316 34700
rect 17368 34688 17374 34740
rect 17586 34688 17592 34740
rect 17644 34688 17650 34740
rect 22021 34700 22508 34728
rect 8110 34620 8116 34672
rect 8168 34660 8174 34672
rect 11793 34663 11851 34669
rect 11793 34660 11805 34663
rect 8168 34632 11805 34660
rect 8168 34620 8174 34632
rect 11793 34629 11805 34632
rect 11839 34660 11851 34663
rect 16390 34660 16396 34672
rect 11839 34632 16396 34660
rect 11839 34629 11851 34632
rect 11793 34623 11851 34629
rect 16390 34620 16396 34632
rect 16448 34620 16454 34672
rect 16758 34620 16764 34672
rect 16816 34660 16822 34672
rect 17221 34663 17279 34669
rect 17221 34660 17233 34663
rect 16816 34632 17233 34660
rect 16816 34620 16822 34632
rect 17221 34629 17233 34632
rect 17267 34660 17279 34663
rect 17604 34660 17632 34688
rect 17267 34632 17632 34660
rect 17267 34629 17279 34632
rect 17221 34623 17279 34629
rect 20990 34620 20996 34672
rect 21048 34620 21054 34672
rect 21266 34669 21272 34672
rect 21209 34663 21272 34669
rect 21209 34629 21221 34663
rect 21255 34629 21272 34663
rect 21209 34623 21272 34629
rect 21266 34620 21272 34623
rect 21324 34620 21330 34672
rect 7883 34564 7972 34592
rect 7883 34561 7895 34564
rect 7837 34555 7895 34561
rect 8202 34552 8208 34604
rect 8260 34592 8266 34604
rect 11698 34601 11704 34604
rect 8297 34595 8355 34601
rect 8297 34592 8309 34595
rect 8260 34564 8309 34592
rect 8260 34552 8266 34564
rect 8297 34561 8309 34564
rect 8343 34561 8355 34595
rect 11696 34592 11704 34601
rect 11659 34564 11704 34592
rect 8297 34555 8355 34561
rect 11696 34555 11704 34564
rect 11698 34552 11704 34555
rect 11756 34552 11762 34604
rect 11885 34595 11943 34601
rect 11885 34561 11897 34595
rect 11931 34592 11943 34595
rect 11974 34592 11980 34604
rect 11931 34564 11980 34592
rect 11931 34561 11943 34564
rect 11885 34555 11943 34561
rect 11974 34552 11980 34564
rect 12032 34552 12038 34604
rect 12068 34595 12126 34601
rect 12068 34561 12080 34595
rect 12114 34561 12126 34595
rect 12068 34555 12126 34561
rect 12161 34595 12219 34601
rect 12161 34561 12173 34595
rect 12207 34592 12219 34595
rect 12250 34592 12256 34604
rect 12207 34564 12256 34592
rect 12207 34561 12219 34564
rect 12161 34555 12219 34561
rect 8389 34527 8447 34533
rect 8389 34493 8401 34527
rect 8435 34493 8447 34527
rect 8389 34487 8447 34493
rect 8573 34527 8631 34533
rect 8573 34493 8585 34527
rect 8619 34524 8631 34527
rect 8846 34524 8852 34536
rect 8619 34496 8852 34524
rect 8619 34493 8631 34496
rect 8573 34487 8631 34493
rect 8404 34456 8432 34487
rect 8846 34484 8852 34496
rect 8904 34484 8910 34536
rect 12084 34524 12112 34555
rect 12250 34552 12256 34564
rect 12308 34552 12314 34604
rect 17126 34592 17132 34604
rect 14016 34564 17132 34592
rect 12084 34496 12434 34524
rect 8662 34456 8668 34468
rect 8404 34428 8668 34456
rect 8662 34416 8668 34428
rect 8720 34456 8726 34468
rect 11790 34456 11796 34468
rect 8720 34428 11796 34456
rect 8720 34416 8726 34428
rect 11790 34416 11796 34428
rect 11848 34416 11854 34468
rect 5350 34348 5356 34400
rect 5408 34388 5414 34400
rect 5445 34391 5503 34397
rect 5445 34388 5457 34391
rect 5408 34360 5457 34388
rect 5408 34348 5414 34360
rect 5445 34357 5457 34360
rect 5491 34357 5503 34391
rect 5445 34351 5503 34357
rect 8846 34348 8852 34400
rect 8904 34388 8910 34400
rect 9858 34388 9864 34400
rect 8904 34360 9864 34388
rect 8904 34348 8910 34360
rect 9858 34348 9864 34360
rect 9916 34348 9922 34400
rect 11514 34348 11520 34400
rect 11572 34348 11578 34400
rect 12406 34388 12434 34496
rect 14016 34468 14044 34564
rect 17126 34552 17132 34564
rect 17184 34552 17190 34604
rect 22021 34601 22049 34700
rect 22094 34620 22100 34672
rect 22152 34660 22158 34672
rect 22189 34663 22247 34669
rect 22189 34660 22201 34663
rect 22152 34632 22201 34660
rect 22152 34620 22158 34632
rect 22189 34629 22201 34632
rect 22235 34629 22247 34663
rect 22480 34660 22508 34700
rect 22554 34688 22560 34740
rect 22612 34728 22618 34740
rect 23014 34728 23020 34740
rect 22612 34700 23020 34728
rect 22612 34688 22618 34700
rect 23014 34688 23020 34700
rect 23072 34728 23078 34740
rect 23750 34728 23756 34740
rect 23072 34700 23428 34728
rect 23072 34688 23078 34700
rect 23198 34660 23204 34672
rect 22480 34632 23204 34660
rect 22189 34623 22247 34629
rect 23198 34620 23204 34632
rect 23256 34620 23262 34672
rect 21913 34595 21971 34601
rect 17236 34564 19334 34592
rect 14918 34484 14924 34536
rect 14976 34524 14982 34536
rect 17236 34524 17264 34564
rect 14976 34496 17264 34524
rect 14976 34484 14982 34496
rect 13998 34416 14004 34468
rect 14056 34416 14062 34468
rect 19306 34456 19334 34564
rect 21913 34561 21925 34595
rect 21959 34561 21971 34595
rect 21913 34555 21971 34561
rect 22006 34595 22064 34601
rect 22006 34561 22018 34595
rect 22052 34561 22064 34595
rect 22006 34555 22064 34561
rect 21928 34524 21956 34555
rect 22278 34552 22284 34604
rect 22336 34552 22342 34604
rect 22378 34595 22436 34601
rect 22378 34561 22390 34595
rect 22424 34592 22436 34595
rect 23106 34592 23112 34604
rect 22424 34564 23112 34592
rect 22424 34561 22436 34564
rect 22378 34555 22436 34561
rect 22296 34524 22324 34552
rect 21376 34496 21956 34524
rect 22021 34496 22324 34524
rect 21376 34465 21404 34496
rect 21361 34459 21419 34465
rect 16500 34428 18092 34456
rect 19306 34428 21312 34456
rect 12526 34388 12532 34400
rect 12406 34360 12532 34388
rect 12526 34348 12532 34360
rect 12584 34388 12590 34400
rect 13170 34388 13176 34400
rect 12584 34360 13176 34388
rect 12584 34348 12590 34360
rect 13170 34348 13176 34360
rect 13228 34388 13234 34400
rect 16500 34388 16528 34428
rect 18064 34400 18092 34428
rect 13228 34360 16528 34388
rect 13228 34348 13234 34360
rect 16850 34348 16856 34400
rect 16908 34348 16914 34400
rect 16942 34348 16948 34400
rect 17000 34348 17006 34400
rect 17034 34348 17040 34400
rect 17092 34348 17098 34400
rect 18046 34348 18052 34400
rect 18104 34348 18110 34400
rect 20622 34348 20628 34400
rect 20680 34388 20686 34400
rect 21177 34391 21235 34397
rect 21177 34388 21189 34391
rect 20680 34360 21189 34388
rect 20680 34348 20686 34360
rect 21177 34357 21189 34360
rect 21223 34357 21235 34391
rect 21284 34388 21312 34428
rect 21361 34425 21373 34459
rect 21407 34425 21419 34459
rect 21361 34419 21419 34425
rect 22021 34388 22049 34496
rect 22393 34456 22421 34555
rect 23106 34552 23112 34564
rect 23164 34552 23170 34604
rect 23216 34524 23244 34620
rect 23400 34601 23428 34700
rect 23492 34700 23756 34728
rect 23492 34604 23520 34700
rect 23750 34688 23756 34700
rect 23808 34688 23814 34740
rect 25314 34688 25320 34740
rect 25372 34728 25378 34740
rect 26694 34728 26700 34740
rect 25372 34700 26700 34728
rect 25372 34688 25378 34700
rect 26694 34688 26700 34700
rect 26752 34688 26758 34740
rect 28810 34688 28816 34740
rect 28868 34688 28874 34740
rect 30926 34688 30932 34740
rect 30984 34688 30990 34740
rect 31205 34731 31263 34737
rect 31205 34697 31217 34731
rect 31251 34728 31263 34731
rect 31386 34728 31392 34740
rect 31251 34700 31392 34728
rect 31251 34697 31263 34700
rect 31205 34691 31263 34697
rect 31386 34688 31392 34700
rect 31444 34688 31450 34740
rect 33318 34728 33324 34740
rect 31726 34700 33324 34728
rect 23569 34663 23627 34669
rect 23569 34629 23581 34663
rect 23615 34660 23627 34663
rect 23615 34632 25912 34660
rect 23615 34629 23627 34632
rect 23569 34623 23627 34629
rect 23385 34595 23443 34601
rect 23385 34561 23397 34595
rect 23431 34561 23443 34595
rect 23385 34555 23443 34561
rect 23474 34552 23480 34604
rect 23532 34552 23538 34604
rect 23661 34595 23719 34601
rect 23661 34561 23673 34595
rect 23707 34561 23719 34595
rect 23661 34555 23719 34561
rect 23753 34595 23811 34601
rect 23753 34561 23765 34595
rect 23799 34592 23811 34595
rect 23842 34592 23848 34604
rect 23799 34564 23848 34592
rect 23799 34561 23811 34564
rect 23753 34555 23811 34561
rect 23676 34524 23704 34555
rect 23842 34552 23848 34564
rect 23900 34552 23906 34604
rect 25884 34592 25912 34632
rect 25958 34620 25964 34672
rect 26016 34660 26022 34672
rect 26142 34660 26148 34672
rect 26016 34632 26148 34660
rect 26016 34620 26022 34632
rect 26142 34620 26148 34632
rect 26200 34620 26206 34672
rect 28534 34620 28540 34672
rect 28592 34620 28598 34672
rect 28828 34660 28856 34688
rect 28644 34632 28856 34660
rect 30944 34660 30972 34688
rect 31726 34660 31754 34700
rect 33318 34688 33324 34700
rect 33376 34688 33382 34740
rect 33502 34688 33508 34740
rect 33560 34728 33566 34740
rect 33689 34731 33747 34737
rect 33689 34728 33701 34731
rect 33560 34700 33701 34728
rect 33560 34688 33566 34700
rect 33689 34697 33701 34700
rect 33735 34697 33747 34731
rect 33689 34691 33747 34697
rect 30944 34632 31754 34660
rect 26418 34592 26424 34604
rect 25884 34564 26424 34592
rect 26418 34552 26424 34564
rect 26476 34552 26482 34604
rect 23216 34496 23704 34524
rect 28552 34524 28580 34620
rect 28644 34601 28672 34632
rect 28629 34595 28687 34601
rect 28629 34561 28641 34595
rect 28675 34561 28687 34595
rect 28629 34555 28687 34561
rect 30024 34524 30052 34578
rect 31570 34552 31576 34604
rect 31628 34592 31634 34604
rect 31628 34564 33272 34592
rect 31628 34552 31634 34564
rect 28552 34496 30052 34524
rect 31662 34484 31668 34536
rect 31720 34484 31726 34536
rect 31757 34527 31815 34533
rect 31757 34493 31769 34527
rect 31803 34493 31815 34527
rect 31757 34487 31815 34493
rect 24946 34456 24952 34468
rect 22112 34428 22421 34456
rect 23032 34428 24952 34456
rect 22112 34400 22140 34428
rect 23032 34400 23060 34428
rect 24946 34416 24952 34428
rect 25004 34456 25010 34468
rect 26418 34456 26424 34468
rect 25004 34428 26424 34456
rect 25004 34416 25010 34428
rect 26418 34416 26424 34428
rect 26476 34416 26482 34468
rect 30834 34416 30840 34468
rect 30892 34456 30898 34468
rect 31294 34456 31300 34468
rect 30892 34428 31300 34456
rect 30892 34416 30898 34428
rect 31294 34416 31300 34428
rect 31352 34456 31358 34468
rect 31772 34456 31800 34487
rect 32766 34484 32772 34536
rect 32824 34524 32830 34536
rect 33244 34533 33272 34564
rect 36906 34552 36912 34604
rect 36964 34592 36970 34604
rect 37553 34595 37611 34601
rect 37553 34592 37565 34595
rect 36964 34564 37565 34592
rect 36964 34552 36970 34564
rect 37553 34561 37565 34564
rect 37599 34561 37611 34595
rect 37553 34555 37611 34561
rect 33045 34527 33103 34533
rect 33045 34524 33057 34527
rect 32824 34496 33057 34524
rect 32824 34484 32830 34496
rect 33045 34493 33057 34496
rect 33091 34493 33103 34527
rect 33045 34487 33103 34493
rect 33229 34527 33287 34533
rect 33229 34493 33241 34527
rect 33275 34524 33287 34527
rect 34146 34524 34152 34536
rect 33275 34496 34152 34524
rect 33275 34493 33287 34496
rect 33229 34487 33287 34493
rect 34146 34484 34152 34496
rect 34204 34484 34210 34536
rect 37829 34527 37887 34533
rect 37829 34493 37841 34527
rect 37875 34524 37887 34527
rect 37918 34524 37924 34536
rect 37875 34496 37924 34524
rect 37875 34493 37887 34496
rect 37829 34487 37887 34493
rect 37918 34484 37924 34496
rect 37976 34484 37982 34536
rect 31352 34428 31800 34456
rect 31352 34416 31358 34428
rect 21284 34360 22049 34388
rect 21177 34351 21235 34357
rect 22094 34348 22100 34400
rect 22152 34348 22158 34400
rect 22278 34348 22284 34400
rect 22336 34388 22342 34400
rect 22557 34391 22615 34397
rect 22557 34388 22569 34391
rect 22336 34360 22569 34388
rect 22336 34348 22342 34360
rect 22557 34357 22569 34360
rect 22603 34357 22615 34391
rect 22557 34351 22615 34357
rect 23014 34348 23020 34400
rect 23072 34348 23078 34400
rect 23750 34348 23756 34400
rect 23808 34388 23814 34400
rect 23937 34391 23995 34397
rect 23937 34388 23949 34391
rect 23808 34360 23949 34388
rect 23808 34348 23814 34360
rect 23937 34357 23949 34360
rect 23983 34357 23995 34391
rect 23937 34351 23995 34357
rect 24762 34348 24768 34400
rect 24820 34388 24826 34400
rect 27246 34388 27252 34400
rect 24820 34360 27252 34388
rect 24820 34348 24826 34360
rect 27246 34348 27252 34360
rect 27304 34348 27310 34400
rect 28074 34348 28080 34400
rect 28132 34388 28138 34400
rect 28886 34391 28944 34397
rect 28886 34388 28898 34391
rect 28132 34360 28898 34388
rect 28132 34348 28138 34360
rect 28886 34357 28898 34360
rect 28932 34357 28944 34391
rect 28886 34351 28944 34357
rect 29638 34348 29644 34400
rect 29696 34388 29702 34400
rect 30377 34391 30435 34397
rect 30377 34388 30389 34391
rect 29696 34360 30389 34388
rect 29696 34348 29702 34360
rect 30377 34357 30389 34360
rect 30423 34388 30435 34391
rect 30558 34388 30564 34400
rect 30423 34360 30564 34388
rect 30423 34357 30435 34360
rect 30377 34351 30435 34357
rect 30558 34348 30564 34360
rect 30616 34348 30622 34400
rect 30650 34348 30656 34400
rect 30708 34388 30714 34400
rect 32784 34388 32812 34484
rect 30708 34360 32812 34388
rect 30708 34348 30714 34360
rect 1104 34298 38272 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38272 34298
rect 1104 34224 38272 34246
rect 14826 34184 14832 34196
rect 14384 34156 14832 34184
rect 14384 34128 14412 34156
rect 14826 34144 14832 34156
rect 14884 34144 14890 34196
rect 15105 34187 15163 34193
rect 15105 34153 15117 34187
rect 15151 34184 15163 34187
rect 16482 34184 16488 34196
rect 15151 34156 16488 34184
rect 15151 34153 15163 34156
rect 15105 34147 15163 34153
rect 16482 34144 16488 34156
rect 16540 34144 16546 34196
rect 16669 34187 16727 34193
rect 16669 34153 16681 34187
rect 16715 34184 16727 34187
rect 16850 34184 16856 34196
rect 16715 34156 16856 34184
rect 16715 34153 16727 34156
rect 16669 34147 16727 34153
rect 16850 34144 16856 34156
rect 16908 34144 16914 34196
rect 16942 34144 16948 34196
rect 17000 34144 17006 34196
rect 17126 34144 17132 34196
rect 17184 34184 17190 34196
rect 17310 34184 17316 34196
rect 17184 34156 17316 34184
rect 17184 34144 17190 34156
rect 17310 34144 17316 34156
rect 17368 34144 17374 34196
rect 17954 34144 17960 34196
rect 18012 34184 18018 34196
rect 18012 34156 26648 34184
rect 18012 34144 18018 34156
rect 11609 34119 11667 34125
rect 11609 34085 11621 34119
rect 11655 34116 11667 34119
rect 14274 34116 14280 34128
rect 11655 34088 14280 34116
rect 11655 34085 11667 34088
rect 11609 34079 11667 34085
rect 14274 34076 14280 34088
rect 14332 34076 14338 34128
rect 14366 34076 14372 34128
rect 14424 34076 14430 34128
rect 14458 34076 14464 34128
rect 14516 34116 14522 34128
rect 15933 34119 15991 34125
rect 14516 34088 15424 34116
rect 14516 34076 14522 34088
rect 15396 34060 15424 34088
rect 15933 34085 15945 34119
rect 15979 34116 15991 34119
rect 16960 34116 16988 34144
rect 17770 34116 17776 34128
rect 15979 34088 16988 34116
rect 17098 34088 17776 34116
rect 15979 34085 15991 34088
rect 15933 34079 15991 34085
rect 5718 34048 5724 34060
rect 4724 34020 5724 34048
rect 4724 33989 4752 34020
rect 5718 34008 5724 34020
rect 5776 34008 5782 34060
rect 9030 34048 9036 34060
rect 8588 34020 9036 34048
rect 4709 33983 4767 33989
rect 4709 33949 4721 33983
rect 4755 33949 4767 33983
rect 4709 33943 4767 33949
rect 4801 33983 4859 33989
rect 4801 33949 4813 33983
rect 4847 33980 4859 33983
rect 4985 33983 5043 33989
rect 4985 33980 4997 33983
rect 4847 33952 4997 33980
rect 4847 33949 4859 33952
rect 4801 33943 4859 33949
rect 4985 33949 4997 33952
rect 5031 33949 5043 33983
rect 4985 33943 5043 33949
rect 6362 33940 6368 33992
rect 6420 33980 6426 33992
rect 6822 33980 6828 33992
rect 6420 33952 6828 33980
rect 6420 33940 6426 33952
rect 6822 33940 6828 33952
rect 6880 33940 6886 33992
rect 7282 33940 7288 33992
rect 7340 33940 7346 33992
rect 8588 33989 8616 34020
rect 9030 34008 9036 34020
rect 9088 34008 9094 34060
rect 12066 34048 12072 34060
rect 9416 34020 12072 34048
rect 8573 33983 8631 33989
rect 8573 33949 8585 33983
rect 8619 33949 8631 33983
rect 8573 33943 8631 33949
rect 5261 33915 5319 33921
rect 5261 33881 5273 33915
rect 5307 33912 5319 33915
rect 5350 33912 5356 33924
rect 5307 33884 5356 33912
rect 5307 33881 5319 33884
rect 5261 33875 5319 33881
rect 5350 33872 5356 33884
rect 5408 33872 5414 33924
rect 9416 33912 9444 34020
rect 12066 34008 12072 34020
rect 12124 34008 12130 34060
rect 13170 34008 13176 34060
rect 13228 34008 13234 34060
rect 13725 34051 13783 34057
rect 13725 34017 13737 34051
rect 13771 34048 13783 34051
rect 14737 34051 14795 34057
rect 14737 34048 14749 34051
rect 13771 34020 14749 34048
rect 13771 34017 13783 34020
rect 13725 34011 13783 34017
rect 14737 34017 14749 34020
rect 14783 34017 14795 34051
rect 14737 34011 14795 34017
rect 15378 34008 15384 34060
rect 15436 34008 15442 34060
rect 16850 34008 16856 34060
rect 16908 34008 16914 34060
rect 17098 34048 17126 34088
rect 17770 34076 17776 34088
rect 17828 34076 17834 34128
rect 19429 34119 19487 34125
rect 18708 34088 19334 34116
rect 18708 34048 18736 34088
rect 17052 34020 17126 34048
rect 17604 34020 18736 34048
rect 19306 34048 19334 34088
rect 19429 34085 19441 34119
rect 19475 34116 19487 34119
rect 19889 34119 19947 34125
rect 19889 34116 19901 34119
rect 19475 34088 19901 34116
rect 19475 34085 19487 34088
rect 19429 34079 19487 34085
rect 19889 34085 19901 34088
rect 19935 34085 19947 34119
rect 19889 34079 19947 34085
rect 20530 34076 20536 34128
rect 20588 34116 20594 34128
rect 26053 34119 26111 34125
rect 20588 34088 25800 34116
rect 20588 34076 20594 34088
rect 19306 34020 20024 34048
rect 9493 33983 9551 33989
rect 9493 33949 9505 33983
rect 9539 33949 9551 33983
rect 9493 33943 9551 33949
rect 6886 33884 9444 33912
rect 9508 33912 9536 33943
rect 9858 33940 9864 33992
rect 9916 33940 9922 33992
rect 11514 33940 11520 33992
rect 11572 33980 11578 33992
rect 11609 33983 11667 33989
rect 11609 33980 11621 33983
rect 11572 33952 11621 33980
rect 11572 33940 11578 33952
rect 11609 33949 11621 33952
rect 11655 33949 11667 33983
rect 11609 33943 11667 33949
rect 11790 33940 11796 33992
rect 11848 33940 11854 33992
rect 11885 33983 11943 33989
rect 11885 33949 11897 33983
rect 11931 33949 11943 33983
rect 11885 33943 11943 33949
rect 9582 33912 9588 33924
rect 9508 33884 9588 33912
rect 6730 33804 6736 33856
rect 6788 33844 6794 33856
rect 6886 33844 6914 33884
rect 9582 33872 9588 33884
rect 9640 33872 9646 33924
rect 11900 33856 11928 33943
rect 13354 33940 13360 33992
rect 13412 33980 13418 33992
rect 13449 33983 13507 33989
rect 13449 33980 13461 33983
rect 13412 33952 13461 33980
rect 13412 33940 13418 33952
rect 13449 33949 13461 33952
rect 13495 33949 13507 33983
rect 13449 33943 13507 33949
rect 14369 33983 14427 33989
rect 14369 33949 14381 33983
rect 14415 33949 14427 33983
rect 14369 33943 14427 33949
rect 14384 33912 14412 33943
rect 14458 33940 14464 33992
rect 14516 33980 14522 33992
rect 14553 33983 14611 33989
rect 14553 33980 14565 33983
rect 14516 33952 14565 33980
rect 14516 33940 14522 33952
rect 14553 33949 14565 33952
rect 14599 33949 14611 33983
rect 14553 33943 14611 33949
rect 14645 33983 14703 33989
rect 14645 33949 14657 33983
rect 14691 33949 14703 33983
rect 14645 33943 14703 33949
rect 14384 33884 14596 33912
rect 14568 33856 14596 33884
rect 14660 33856 14688 33943
rect 16022 33940 16028 33992
rect 16080 33940 16086 33992
rect 16206 33940 16212 33992
rect 16264 33940 16270 33992
rect 16298 33940 16304 33992
rect 16356 33940 16362 33992
rect 16390 33940 16396 33992
rect 16448 33940 16454 33992
rect 17052 33989 17080 34020
rect 17037 33983 17095 33989
rect 17037 33949 17049 33983
rect 17083 33949 17095 33983
rect 17037 33943 17095 33949
rect 17126 33940 17132 33992
rect 17184 33980 17190 33992
rect 17221 33983 17279 33989
rect 17221 33980 17233 33983
rect 17184 33952 17233 33980
rect 17184 33940 17190 33952
rect 17221 33949 17233 33952
rect 17267 33949 17279 33983
rect 17221 33943 17279 33949
rect 17310 33940 17316 33992
rect 17368 33940 17374 33992
rect 17405 33983 17463 33989
rect 17405 33949 17417 33983
rect 17451 33980 17463 33983
rect 17604 33980 17632 34020
rect 17451 33952 17632 33980
rect 17451 33949 17463 33952
rect 17405 33943 17463 33949
rect 17678 33940 17684 33992
rect 17736 33940 17742 33992
rect 17774 33983 17832 33989
rect 17774 33949 17786 33983
rect 17820 33949 17832 33983
rect 17774 33943 17832 33949
rect 18146 33983 18204 33989
rect 18146 33949 18158 33983
rect 18192 33949 18204 33983
rect 18146 33943 18204 33949
rect 15565 33915 15623 33921
rect 15565 33881 15577 33915
rect 15611 33912 15623 33915
rect 17328 33912 17356 33940
rect 17789 33912 17817 33943
rect 15611 33884 16620 33912
rect 17328 33884 17817 33912
rect 15611 33881 15623 33884
rect 15565 33875 15623 33881
rect 6788 33816 6914 33844
rect 6788 33804 6794 33816
rect 7190 33804 7196 33856
rect 7248 33804 7254 33856
rect 8662 33804 8668 33856
rect 8720 33804 8726 33856
rect 8938 33804 8944 33856
rect 8996 33804 9002 33856
rect 9398 33804 9404 33856
rect 9456 33844 9462 33856
rect 9677 33847 9735 33853
rect 9677 33844 9689 33847
rect 9456 33816 9689 33844
rect 9456 33804 9462 33816
rect 9677 33813 9689 33816
rect 9723 33813 9735 33847
rect 9677 33807 9735 33813
rect 11882 33804 11888 33856
rect 11940 33804 11946 33856
rect 13262 33804 13268 33856
rect 13320 33844 13326 33856
rect 13357 33847 13415 33853
rect 13357 33844 13369 33847
rect 13320 33816 13369 33844
rect 13320 33804 13326 33816
rect 13357 33813 13369 33816
rect 13403 33813 13415 33847
rect 13357 33807 13415 33813
rect 13541 33847 13599 33853
rect 13541 33813 13553 33847
rect 13587 33844 13599 33847
rect 13722 33844 13728 33856
rect 13587 33816 13728 33844
rect 13587 33813 13599 33816
rect 13541 33807 13599 33813
rect 13722 33804 13728 33816
rect 13780 33804 13786 33856
rect 14550 33804 14556 33856
rect 14608 33804 14614 33856
rect 14642 33804 14648 33856
rect 14700 33804 14706 33856
rect 15654 33804 15660 33856
rect 15712 33804 15718 33856
rect 15749 33847 15807 33853
rect 15749 33813 15761 33847
rect 15795 33844 15807 33847
rect 16022 33844 16028 33856
rect 15795 33816 16028 33844
rect 15795 33813 15807 33816
rect 15749 33807 15807 33813
rect 16022 33804 16028 33816
rect 16080 33844 16086 33856
rect 16390 33844 16396 33856
rect 16080 33816 16396 33844
rect 16080 33804 16086 33816
rect 16390 33804 16396 33816
rect 16448 33804 16454 33856
rect 16592 33844 16620 33884
rect 17954 33872 17960 33924
rect 18012 33872 18018 33924
rect 18046 33872 18052 33924
rect 18104 33872 18110 33924
rect 16942 33844 16948 33856
rect 16592 33816 16948 33844
rect 16942 33804 16948 33816
rect 17000 33804 17006 33856
rect 17131 33853 17137 33856
rect 17129 33807 17137 33853
rect 17189 33844 17195 33856
rect 17189 33816 17229 33844
rect 17131 33804 17137 33807
rect 17189 33804 17195 33816
rect 17310 33804 17316 33856
rect 17368 33844 17374 33856
rect 18161 33844 18189 33943
rect 18414 33940 18420 33992
rect 18472 33940 18478 33992
rect 18693 33983 18751 33989
rect 18693 33980 18705 33983
rect 18524 33952 18705 33980
rect 18230 33872 18236 33924
rect 18288 33912 18294 33924
rect 18524 33912 18552 33952
rect 18693 33949 18705 33952
rect 18739 33949 18751 33983
rect 18693 33943 18751 33949
rect 18288 33884 18552 33912
rect 18288 33872 18294 33884
rect 18598 33872 18604 33924
rect 18656 33872 18662 33924
rect 18708 33912 18736 33943
rect 18782 33940 18788 33992
rect 18840 33940 18846 33992
rect 19242 33940 19248 33992
rect 19300 33940 19306 33992
rect 19521 33983 19579 33989
rect 19521 33980 19533 33983
rect 19352 33952 19533 33980
rect 19058 33912 19064 33924
rect 18708 33884 19064 33912
rect 19058 33872 19064 33884
rect 19116 33872 19122 33924
rect 17368 33816 18189 33844
rect 17368 33804 17374 33816
rect 18322 33804 18328 33856
rect 18380 33804 18386 33856
rect 18969 33847 19027 33853
rect 18969 33813 18981 33847
rect 19015 33844 19027 33847
rect 19352 33844 19380 33952
rect 19521 33949 19533 33952
rect 19567 33949 19579 33983
rect 19521 33943 19579 33949
rect 19996 33912 20024 34020
rect 20088 34020 21772 34048
rect 20088 33989 20116 34020
rect 21744 33992 21772 34020
rect 22204 34020 25728 34048
rect 20073 33983 20131 33989
rect 20073 33949 20085 33983
rect 20119 33949 20131 33983
rect 20073 33943 20131 33949
rect 20254 33940 20260 33992
rect 20312 33940 20318 33992
rect 20441 33983 20499 33989
rect 20441 33949 20453 33983
rect 20487 33980 20499 33983
rect 20530 33980 20536 33992
rect 20487 33952 20536 33980
rect 20487 33949 20499 33952
rect 20441 33943 20499 33949
rect 20530 33940 20536 33952
rect 20588 33940 20594 33992
rect 20622 33940 20628 33992
rect 20680 33980 20686 33992
rect 20809 33983 20867 33989
rect 20809 33980 20821 33983
rect 20680 33952 20821 33980
rect 20680 33940 20686 33952
rect 20809 33949 20821 33952
rect 20855 33949 20867 33983
rect 20809 33943 20867 33949
rect 21726 33940 21732 33992
rect 21784 33940 21790 33992
rect 21910 33940 21916 33992
rect 21968 33940 21974 33992
rect 22094 33940 22100 33992
rect 22152 33940 22158 33992
rect 20165 33915 20223 33921
rect 20165 33912 20177 33915
rect 19996 33884 20177 33912
rect 20165 33881 20177 33884
rect 20211 33912 20223 33915
rect 22204 33912 22232 34020
rect 22278 33940 22284 33992
rect 22336 33940 22342 33992
rect 22462 33940 22468 33992
rect 22520 33980 22526 33992
rect 22557 33983 22615 33989
rect 22557 33980 22569 33983
rect 22520 33952 22569 33980
rect 22520 33940 22526 33952
rect 22557 33949 22569 33952
rect 22603 33949 22615 33983
rect 22557 33943 22615 33949
rect 22649 33983 22707 33989
rect 22649 33949 22661 33983
rect 22695 33949 22707 33983
rect 22649 33943 22707 33949
rect 22833 33983 22891 33989
rect 22833 33949 22845 33983
rect 22879 33949 22891 33983
rect 22833 33943 22891 33949
rect 22925 33983 22983 33989
rect 22925 33949 22937 33983
rect 22971 33949 22983 33983
rect 22925 33943 22983 33949
rect 20211 33884 22232 33912
rect 22296 33912 22324 33940
rect 22664 33912 22692 33943
rect 22296 33884 22692 33912
rect 20211 33881 20223 33884
rect 20165 33875 20223 33881
rect 19015 33816 19380 33844
rect 19521 33847 19579 33853
rect 19015 33813 19027 33816
rect 18969 33807 19027 33813
rect 19521 33813 19533 33847
rect 19567 33844 19579 33847
rect 20346 33844 20352 33856
rect 19567 33816 20352 33844
rect 19567 33813 19579 33816
rect 19521 33807 19579 33813
rect 20346 33804 20352 33816
rect 20404 33804 20410 33856
rect 21726 33804 21732 33856
rect 21784 33844 21790 33856
rect 22462 33844 22468 33856
rect 21784 33816 22468 33844
rect 21784 33804 21790 33816
rect 22462 33804 22468 33816
rect 22520 33804 22526 33856
rect 22554 33804 22560 33856
rect 22612 33844 22618 33856
rect 22848 33844 22876 33943
rect 22612 33816 22876 33844
rect 22940 33844 22968 33943
rect 23198 33940 23204 33992
rect 23256 33940 23262 33992
rect 23294 33983 23352 33989
rect 23294 33949 23306 33983
rect 23340 33949 23352 33983
rect 23294 33943 23352 33949
rect 23308 33912 23336 33943
rect 23474 33940 23480 33992
rect 23532 33940 23538 33992
rect 23566 33940 23572 33992
rect 23624 33940 23630 33992
rect 23707 33983 23765 33989
rect 23707 33949 23719 33983
rect 23753 33980 23765 33983
rect 24210 33980 24216 33992
rect 23753 33952 24216 33980
rect 23753 33949 23765 33952
rect 23707 33943 23765 33949
rect 24210 33940 24216 33952
rect 24268 33980 24274 33992
rect 24762 33980 24768 33992
rect 24268 33952 24768 33980
rect 24268 33940 24274 33952
rect 24762 33940 24768 33952
rect 24820 33940 24826 33992
rect 25406 33940 25412 33992
rect 25464 33980 25470 33992
rect 25700 33989 25728 34020
rect 25593 33983 25651 33989
rect 25593 33980 25605 33983
rect 25464 33952 25605 33980
rect 25464 33940 25470 33952
rect 25593 33949 25605 33952
rect 25639 33949 25651 33983
rect 25593 33943 25651 33949
rect 25685 33983 25743 33989
rect 25685 33949 25697 33983
rect 25731 33949 25743 33983
rect 25685 33943 25743 33949
rect 24026 33912 24032 33924
rect 23308 33884 24032 33912
rect 24026 33872 24032 33884
rect 24084 33872 24090 33924
rect 25608 33912 25636 33943
rect 24504 33884 25636 33912
rect 24504 33856 24532 33884
rect 23014 33844 23020 33856
rect 22940 33816 23020 33844
rect 22612 33804 22618 33816
rect 23014 33804 23020 33816
rect 23072 33804 23078 33856
rect 23106 33804 23112 33856
rect 23164 33804 23170 33856
rect 23842 33804 23848 33856
rect 23900 33804 23906 33856
rect 24486 33804 24492 33856
rect 24544 33804 24550 33856
rect 25406 33804 25412 33856
rect 25464 33804 25470 33856
rect 25700 33844 25728 33943
rect 25772 33912 25800 34088
rect 26053 34085 26065 34119
rect 26099 34085 26111 34119
rect 26053 34079 26111 34085
rect 26620 34116 26648 34156
rect 28074 34144 28080 34196
rect 28132 34144 28138 34196
rect 30834 34184 30840 34196
rect 28368 34156 30840 34184
rect 28368 34116 28396 34156
rect 30834 34144 30840 34156
rect 30892 34144 30898 34196
rect 26620 34088 28396 34116
rect 26068 34048 26096 34079
rect 25884 34020 26096 34048
rect 25884 33989 25912 34020
rect 25869 33983 25927 33989
rect 25869 33949 25881 33983
rect 25915 33949 25927 33983
rect 25869 33943 25927 33949
rect 25958 33940 25964 33992
rect 26016 33940 26022 33992
rect 26142 33940 26148 33992
rect 26200 33980 26206 33992
rect 26620 33989 26648 34088
rect 28442 34076 28448 34128
rect 28500 34076 28506 34128
rect 28644 34088 29777 34116
rect 28644 34048 28672 34088
rect 29089 34051 29147 34057
rect 29089 34048 29101 34051
rect 26712 34020 28672 34048
rect 28966 34020 29101 34048
rect 26237 33983 26295 33989
rect 26237 33980 26249 33983
rect 26200 33952 26249 33980
rect 26200 33940 26206 33952
rect 26237 33949 26249 33952
rect 26283 33949 26295 33983
rect 26237 33943 26295 33949
rect 26329 33983 26387 33989
rect 26329 33949 26341 33983
rect 26375 33980 26387 33983
rect 26605 33983 26663 33989
rect 26375 33952 26556 33980
rect 26375 33949 26387 33952
rect 26329 33943 26387 33949
rect 26344 33912 26372 33943
rect 25772 33884 26372 33912
rect 26418 33872 26424 33924
rect 26476 33872 26482 33924
rect 26528 33912 26556 33952
rect 26605 33949 26617 33983
rect 26651 33949 26663 33983
rect 26605 33943 26663 33949
rect 26712 33912 26740 34020
rect 26970 33940 26976 33992
rect 27028 33980 27034 33992
rect 27249 33983 27307 33989
rect 27249 33980 27261 33983
rect 27028 33952 27261 33980
rect 27028 33940 27034 33952
rect 27249 33949 27261 33952
rect 27295 33949 27307 33983
rect 27249 33943 27307 33949
rect 27893 33983 27951 33989
rect 27893 33949 27905 33983
rect 27939 33980 27951 33983
rect 28442 33980 28448 33992
rect 27939 33952 28448 33980
rect 27939 33949 27951 33952
rect 27893 33943 27951 33949
rect 28442 33940 28448 33952
rect 28500 33940 28506 33992
rect 28626 33940 28632 33992
rect 28684 33980 28690 33992
rect 28966 33980 28994 34020
rect 29089 34017 29101 34020
rect 29135 34017 29147 34051
rect 29089 34011 29147 34017
rect 28684 33952 28994 33980
rect 28684 33940 28690 33952
rect 28905 33915 28963 33921
rect 28905 33912 28917 33915
rect 26528 33884 26740 33912
rect 26804 33884 28917 33912
rect 26804 33844 26832 33884
rect 28905 33881 28917 33884
rect 28951 33881 28963 33915
rect 28905 33875 28963 33881
rect 25700 33816 26832 33844
rect 27154 33804 27160 33856
rect 27212 33804 27218 33856
rect 28166 33804 28172 33856
rect 28224 33844 28230 33856
rect 28810 33844 28816 33856
rect 28224 33816 28816 33844
rect 28224 33804 28230 33816
rect 28810 33804 28816 33816
rect 28868 33804 28874 33856
rect 28920 33844 28948 33875
rect 29638 33844 29644 33856
rect 28920 33816 29644 33844
rect 29638 33804 29644 33816
rect 29696 33804 29702 33856
rect 29749 33844 29777 34088
rect 29914 34076 29920 34128
rect 29972 34116 29978 34128
rect 31113 34119 31171 34125
rect 29972 34088 30972 34116
rect 29972 34076 29978 34088
rect 29822 33940 29828 33992
rect 29880 33940 29886 33992
rect 30466 33940 30472 33992
rect 30524 33940 30530 33992
rect 30558 33940 30564 33992
rect 30616 33980 30622 33992
rect 30616 33952 30661 33980
rect 30616 33940 30622 33952
rect 30834 33940 30840 33992
rect 30892 33940 30898 33992
rect 30944 33989 30972 34088
rect 31113 34085 31125 34119
rect 31159 34116 31171 34119
rect 34057 34119 34115 34125
rect 31159 34088 31754 34116
rect 31159 34085 31171 34088
rect 31113 34079 31171 34085
rect 31726 34048 31754 34088
rect 34057 34085 34069 34119
rect 34103 34085 34115 34119
rect 34057 34079 34115 34085
rect 34072 34048 34100 34079
rect 34977 34051 35035 34057
rect 34977 34048 34989 34051
rect 31726 34020 31800 34048
rect 34072 34020 34989 34048
rect 30934 33983 30992 33989
rect 30934 33949 30946 33983
rect 30980 33949 30992 33983
rect 30934 33943 30992 33949
rect 31478 33940 31484 33992
rect 31536 33940 31542 33992
rect 31772 33989 31800 34020
rect 34977 34017 34989 34020
rect 35023 34017 35035 34051
rect 34977 34011 35035 34017
rect 31757 33983 31815 33989
rect 31757 33949 31769 33983
rect 31803 33949 31815 33983
rect 31757 33943 31815 33949
rect 33870 33940 33876 33992
rect 33928 33940 33934 33992
rect 34330 33940 34336 33992
rect 34388 33940 34394 33992
rect 34425 33983 34483 33989
rect 34425 33949 34437 33983
rect 34471 33980 34483 33983
rect 34701 33983 34759 33989
rect 34701 33980 34713 33983
rect 34471 33952 34713 33980
rect 34471 33949 34483 33952
rect 34425 33943 34483 33949
rect 34701 33949 34713 33952
rect 34747 33949 34759 33983
rect 34701 33943 34759 33949
rect 29840 33912 29868 33940
rect 30745 33915 30803 33921
rect 30745 33912 30757 33915
rect 29840 33884 30757 33912
rect 30745 33881 30757 33884
rect 30791 33881 30803 33915
rect 30745 33875 30803 33881
rect 34256 33884 35466 33912
rect 31573 33847 31631 33853
rect 31573 33844 31585 33847
rect 29749 33816 31585 33844
rect 31573 33813 31585 33816
rect 31619 33844 31631 33847
rect 31662 33844 31668 33856
rect 31619 33816 31668 33844
rect 31619 33813 31631 33816
rect 31573 33807 31631 33813
rect 31662 33804 31668 33816
rect 31720 33804 31726 33856
rect 31941 33847 31999 33853
rect 31941 33813 31953 33847
rect 31987 33844 31999 33847
rect 32214 33844 32220 33856
rect 31987 33816 32220 33844
rect 31987 33813 31999 33816
rect 31941 33807 31999 33813
rect 32214 33804 32220 33816
rect 32272 33804 32278 33856
rect 33318 33804 33324 33856
rect 33376 33844 33382 33856
rect 34256 33844 34284 33884
rect 33376 33816 34284 33844
rect 35360 33844 35388 33884
rect 36262 33872 36268 33924
rect 36320 33912 36326 33924
rect 36725 33915 36783 33921
rect 36725 33912 36737 33915
rect 36320 33884 36737 33912
rect 36320 33872 36326 33884
rect 36725 33881 36737 33884
rect 36771 33881 36783 33915
rect 36725 33875 36783 33881
rect 35986 33844 35992 33856
rect 35360 33816 35992 33844
rect 33376 33804 33382 33816
rect 35986 33804 35992 33816
rect 36044 33804 36050 33856
rect 1104 33754 38272 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38272 33754
rect 1104 33680 38272 33702
rect 5445 33643 5503 33649
rect 5445 33609 5457 33643
rect 5491 33640 5503 33643
rect 5534 33640 5540 33652
rect 5491 33612 5540 33640
rect 5491 33609 5503 33612
rect 5445 33603 5503 33609
rect 5534 33600 5540 33612
rect 5592 33600 5598 33652
rect 5813 33643 5871 33649
rect 5813 33609 5825 33643
rect 5859 33640 5871 33643
rect 6730 33640 6736 33652
rect 5859 33612 6736 33640
rect 5859 33609 5871 33612
rect 5813 33603 5871 33609
rect 6730 33600 6736 33612
rect 6788 33600 6794 33652
rect 7190 33600 7196 33652
rect 7248 33600 7254 33652
rect 8662 33600 8668 33652
rect 8720 33600 8726 33652
rect 9398 33640 9404 33652
rect 9232 33612 9404 33640
rect 7208 33572 7236 33600
rect 7024 33544 7236 33572
rect 7024 33513 7052 33544
rect 7009 33507 7067 33513
rect 7009 33473 7021 33507
rect 7055 33473 7067 33507
rect 7009 33467 7067 33473
rect 8294 33464 8300 33516
rect 8352 33504 8358 33516
rect 8680 33504 8708 33600
rect 9232 33581 9260 33612
rect 9398 33600 9404 33612
rect 9456 33600 9462 33652
rect 13354 33600 13360 33652
rect 13412 33600 13418 33652
rect 13906 33600 13912 33652
rect 13964 33640 13970 33652
rect 14369 33643 14427 33649
rect 14369 33640 14381 33643
rect 13964 33612 14381 33640
rect 13964 33600 13970 33612
rect 14369 33609 14381 33612
rect 14415 33609 14427 33643
rect 14369 33603 14427 33609
rect 14553 33643 14611 33649
rect 14553 33609 14565 33643
rect 14599 33640 14611 33643
rect 14642 33640 14648 33652
rect 14599 33612 14648 33640
rect 14599 33609 14611 33612
rect 14553 33603 14611 33609
rect 14642 33600 14648 33612
rect 14700 33600 14706 33652
rect 16666 33600 16672 33652
rect 16724 33640 16730 33652
rect 17310 33640 17316 33652
rect 16724 33612 17316 33640
rect 16724 33600 16730 33612
rect 17310 33600 17316 33612
rect 17368 33600 17374 33652
rect 17589 33643 17647 33649
rect 17589 33609 17601 33643
rect 17635 33640 17647 33643
rect 17678 33640 17684 33652
rect 17635 33612 17684 33640
rect 17635 33609 17647 33612
rect 17589 33603 17647 33609
rect 17678 33600 17684 33612
rect 17736 33600 17742 33652
rect 19334 33600 19340 33652
rect 19392 33640 19398 33652
rect 19392 33612 19932 33640
rect 19392 33600 19398 33612
rect 9217 33575 9275 33581
rect 9217 33541 9229 33575
rect 9263 33541 9275 33575
rect 9217 33535 9275 33541
rect 11790 33532 11796 33584
rect 11848 33572 11854 33584
rect 13372 33572 13400 33600
rect 14277 33575 14335 33581
rect 14277 33572 14289 33575
rect 11848 33544 13216 33572
rect 13372 33544 14289 33572
rect 11848 33532 11854 33544
rect 8941 33507 8999 33513
rect 8941 33504 8953 33507
rect 8352 33476 8418 33504
rect 8680 33476 8953 33504
rect 8352 33464 8358 33476
rect 8941 33473 8953 33476
rect 8987 33473 8999 33507
rect 8941 33467 8999 33473
rect 10318 33464 10324 33516
rect 10376 33464 10382 33516
rect 5902 33396 5908 33448
rect 5960 33396 5966 33448
rect 6089 33439 6147 33445
rect 6089 33405 6101 33439
rect 6135 33436 6147 33439
rect 6135 33408 6914 33436
rect 6135 33405 6147 33408
rect 6089 33399 6147 33405
rect 6886 33300 6914 33408
rect 7282 33396 7288 33448
rect 7340 33396 7346 33448
rect 8757 33439 8815 33445
rect 8757 33405 8769 33439
rect 8803 33436 8815 33439
rect 9582 33436 9588 33448
rect 8803 33408 9588 33436
rect 8803 33405 8815 33408
rect 8757 33399 8815 33405
rect 9582 33396 9588 33408
rect 9640 33436 9646 33448
rect 13188 33436 13216 33544
rect 14277 33541 14289 33544
rect 14323 33541 14335 33575
rect 14277 33535 14335 33541
rect 16482 33532 16488 33584
rect 16540 33572 16546 33584
rect 17221 33575 17279 33581
rect 17221 33572 17233 33575
rect 16540 33544 17233 33572
rect 16540 33532 16546 33544
rect 17221 33541 17233 33544
rect 17267 33541 17279 33575
rect 17221 33535 17279 33541
rect 17451 33541 17509 33547
rect 13262 33464 13268 33516
rect 13320 33504 13326 33516
rect 13538 33504 13544 33516
rect 13320 33476 13544 33504
rect 13320 33464 13326 33476
rect 13538 33464 13544 33476
rect 13596 33504 13602 33516
rect 14185 33507 14243 33513
rect 14185 33504 14197 33507
rect 13596 33476 14197 33504
rect 13596 33464 13602 33476
rect 14185 33473 14197 33476
rect 14231 33473 14243 33507
rect 14185 33467 14243 33473
rect 13998 33436 14004 33448
rect 9640 33408 12296 33436
rect 13188 33408 14004 33436
rect 9640 33396 9646 33408
rect 12268 33368 12296 33408
rect 13998 33396 14004 33408
rect 14056 33396 14062 33448
rect 17236 33436 17264 33535
rect 17451 33507 17463 33541
rect 17497 33507 17509 33541
rect 17451 33504 17509 33507
rect 17770 33504 17776 33516
rect 17451 33501 17776 33504
rect 17466 33476 17776 33501
rect 17236 33408 17540 33436
rect 15746 33368 15752 33380
rect 12268 33340 15752 33368
rect 15746 33328 15752 33340
rect 15804 33328 15810 33380
rect 7466 33300 7472 33312
rect 6886 33272 7472 33300
rect 7466 33260 7472 33272
rect 7524 33260 7530 33312
rect 10594 33260 10600 33312
rect 10652 33300 10658 33312
rect 10689 33303 10747 33309
rect 10689 33300 10701 33303
rect 10652 33272 10701 33300
rect 10652 33260 10658 33272
rect 10689 33269 10701 33272
rect 10735 33300 10747 33303
rect 11790 33300 11796 33312
rect 10735 33272 11796 33300
rect 10735 33269 10747 33272
rect 10689 33263 10747 33269
rect 11790 33260 11796 33272
rect 11848 33260 11854 33312
rect 16206 33260 16212 33312
rect 16264 33300 16270 33312
rect 17405 33303 17463 33309
rect 17405 33300 17417 33303
rect 16264 33272 17417 33300
rect 16264 33260 16270 33272
rect 17405 33269 17417 33272
rect 17451 33269 17463 33303
rect 17512 33300 17540 33408
rect 17604 33380 17632 33476
rect 17770 33464 17776 33476
rect 17828 33464 17834 33516
rect 19702 33513 19708 33516
rect 19696 33467 19708 33513
rect 19702 33464 19708 33467
rect 19760 33464 19766 33516
rect 19904 33513 19932 33612
rect 20254 33600 20260 33652
rect 20312 33640 20318 33652
rect 20312 33612 20944 33640
rect 20312 33600 20318 33612
rect 20809 33575 20867 33581
rect 20809 33572 20821 33575
rect 20272 33544 20821 33572
rect 20272 33513 20300 33544
rect 20809 33541 20821 33544
rect 20855 33541 20867 33575
rect 20916 33572 20944 33612
rect 21082 33600 21088 33652
rect 21140 33600 21146 33652
rect 21266 33600 21272 33652
rect 21324 33640 21330 33652
rect 21910 33640 21916 33652
rect 21324 33612 21916 33640
rect 21324 33600 21330 33612
rect 21910 33600 21916 33612
rect 21968 33600 21974 33652
rect 22462 33600 22468 33652
rect 22520 33640 22526 33652
rect 22646 33640 22652 33652
rect 22520 33612 22652 33640
rect 22520 33600 22526 33612
rect 22646 33600 22652 33612
rect 22704 33600 22710 33652
rect 22830 33600 22836 33652
rect 22888 33640 22894 33652
rect 23014 33640 23020 33652
rect 22888 33612 23020 33640
rect 22888 33600 22894 33612
rect 23014 33600 23020 33612
rect 23072 33600 23078 33652
rect 27154 33600 27160 33652
rect 27212 33600 27218 33652
rect 27338 33600 27344 33652
rect 27396 33640 27402 33652
rect 27396 33612 31754 33640
rect 27396 33600 27402 33612
rect 20916 33544 21404 33572
rect 20809 33535 20867 33541
rect 19889 33507 19947 33513
rect 19889 33473 19901 33507
rect 19935 33473 19947 33507
rect 19889 33467 19947 33473
rect 20257 33507 20315 33513
rect 20257 33473 20269 33507
rect 20303 33473 20315 33507
rect 20257 33467 20315 33473
rect 20346 33464 20352 33516
rect 20404 33464 20410 33516
rect 20622 33464 20628 33516
rect 20680 33464 20686 33516
rect 20717 33507 20775 33513
rect 20717 33473 20729 33507
rect 20763 33504 20775 33507
rect 20901 33507 20959 33513
rect 20763 33476 20852 33504
rect 20763 33473 20775 33476
rect 20717 33467 20775 33473
rect 19058 33396 19064 33448
rect 19116 33396 19122 33448
rect 19610 33396 19616 33448
rect 19668 33436 19674 33448
rect 20640 33436 20668 33464
rect 20824 33448 20852 33476
rect 20901 33473 20913 33507
rect 20947 33473 20959 33507
rect 21376 33504 21404 33544
rect 21450 33532 21456 33584
rect 21508 33532 21514 33584
rect 23290 33572 23296 33584
rect 21560 33544 23296 33572
rect 21560 33504 21588 33544
rect 23290 33532 23296 33544
rect 23348 33532 23354 33584
rect 25225 33575 25283 33581
rect 23676 33544 23980 33572
rect 21376 33476 21588 33504
rect 20901 33467 20959 33473
rect 19668 33408 20668 33436
rect 19668 33396 19674 33408
rect 20806 33396 20812 33448
rect 20864 33396 20870 33448
rect 20916 33436 20944 33467
rect 21818 33464 21824 33516
rect 21876 33464 21882 33516
rect 22005 33507 22063 33513
rect 22005 33504 22017 33507
rect 21928 33476 22017 33504
rect 21928 33436 21956 33476
rect 22005 33473 22017 33476
rect 22051 33504 22063 33507
rect 23676 33504 23704 33544
rect 22051 33476 23704 33504
rect 22051 33473 22063 33476
rect 22005 33467 22063 33473
rect 23750 33464 23756 33516
rect 23808 33464 23814 33516
rect 23842 33464 23848 33516
rect 23900 33464 23906 33516
rect 23952 33504 23980 33544
rect 25225 33541 25237 33575
rect 25271 33572 25283 33575
rect 25314 33572 25320 33584
rect 25271 33544 25320 33572
rect 25271 33541 25283 33544
rect 25225 33535 25283 33541
rect 25314 33532 25320 33544
rect 25372 33532 25378 33584
rect 27172 33572 27200 33600
rect 28534 33572 28540 33584
rect 26988 33544 27200 33572
rect 28474 33544 28540 33572
rect 23952 33476 26556 33504
rect 20916 33408 21956 33436
rect 23474 33396 23480 33448
rect 23532 33396 23538 33448
rect 23569 33439 23627 33445
rect 23569 33405 23581 33439
rect 23615 33436 23627 33439
rect 23934 33436 23940 33448
rect 23615 33408 23940 33436
rect 23615 33405 23627 33408
rect 23569 33399 23627 33405
rect 23934 33396 23940 33408
rect 23992 33396 23998 33448
rect 25406 33396 25412 33448
rect 25464 33396 25470 33448
rect 17586 33328 17592 33380
rect 17644 33328 17650 33380
rect 18138 33328 18144 33380
rect 18196 33368 18202 33380
rect 19886 33368 19892 33380
rect 18196 33340 19892 33368
rect 18196 33328 18202 33340
rect 19886 33328 19892 33340
rect 19944 33328 19950 33380
rect 19978 33328 19984 33380
rect 20036 33368 20042 33380
rect 21821 33371 21879 33377
rect 21821 33368 21833 33371
rect 20036 33340 21833 33368
rect 20036 33328 20042 33340
rect 21821 33337 21833 33340
rect 21867 33368 21879 33371
rect 24857 33371 24915 33377
rect 24857 33368 24869 33371
rect 21867 33340 24869 33368
rect 21867 33337 21879 33340
rect 21821 33331 21879 33337
rect 24857 33337 24869 33340
rect 24903 33337 24915 33371
rect 25424 33368 25452 33396
rect 24857 33331 24915 33337
rect 25240 33340 25452 33368
rect 18414 33300 18420 33312
rect 17512 33272 18420 33300
rect 17405 33263 17463 33269
rect 18414 33260 18420 33272
rect 18472 33260 18478 33312
rect 19426 33260 19432 33312
rect 19484 33300 19490 33312
rect 20530 33300 20536 33312
rect 19484 33272 20536 33300
rect 19484 33260 19490 33272
rect 20530 33260 20536 33272
rect 20588 33260 20594 33312
rect 21269 33303 21327 33309
rect 21269 33269 21281 33303
rect 21315 33300 21327 33303
rect 21450 33300 21456 33312
rect 21315 33272 21456 33300
rect 21315 33269 21327 33272
rect 21269 33263 21327 33269
rect 21450 33260 21456 33272
rect 21508 33260 21514 33312
rect 22094 33260 22100 33312
rect 22152 33300 22158 33312
rect 23842 33300 23848 33312
rect 22152 33272 23848 33300
rect 22152 33260 22158 33272
rect 23842 33260 23848 33272
rect 23900 33260 23906 33312
rect 24026 33260 24032 33312
rect 24084 33260 24090 33312
rect 25240 33309 25268 33340
rect 25225 33303 25283 33309
rect 25225 33269 25237 33303
rect 25271 33269 25283 33303
rect 25225 33263 25283 33269
rect 25406 33260 25412 33312
rect 25464 33260 25470 33312
rect 26528 33300 26556 33476
rect 26602 33464 26608 33516
rect 26660 33464 26666 33516
rect 26988 33513 27016 33544
rect 28534 33532 28540 33544
rect 28592 33532 28598 33584
rect 28810 33532 28816 33584
rect 28868 33572 28874 33584
rect 31570 33572 31576 33584
rect 28868 33544 31576 33572
rect 28868 33532 28874 33544
rect 31570 33532 31576 33544
rect 31628 33532 31634 33584
rect 31726 33572 31754 33612
rect 33134 33600 33140 33652
rect 33192 33640 33198 33652
rect 33321 33643 33379 33649
rect 33321 33640 33333 33643
rect 33192 33612 33333 33640
rect 33192 33600 33198 33612
rect 33321 33609 33333 33612
rect 33367 33609 33379 33643
rect 33321 33603 33379 33609
rect 33781 33643 33839 33649
rect 33781 33609 33793 33643
rect 33827 33640 33839 33643
rect 33870 33640 33876 33652
rect 33827 33612 33876 33640
rect 33827 33609 33839 33612
rect 33781 33603 33839 33609
rect 33870 33600 33876 33612
rect 33928 33600 33934 33652
rect 34146 33600 34152 33652
rect 34204 33600 34210 33652
rect 34609 33643 34667 33649
rect 34609 33609 34621 33643
rect 34655 33609 34667 33643
rect 34609 33603 34667 33609
rect 31726 33544 33456 33572
rect 26973 33507 27031 33513
rect 26973 33473 26985 33507
rect 27019 33473 27031 33507
rect 28552 33504 28580 33532
rect 29178 33504 29184 33516
rect 28552 33476 29184 33504
rect 26973 33467 27031 33473
rect 29178 33464 29184 33476
rect 29236 33504 29242 33516
rect 33318 33504 33324 33516
rect 29236 33476 33324 33504
rect 29236 33464 29242 33476
rect 33318 33464 33324 33476
rect 33376 33464 33382 33516
rect 33428 33513 33456 33544
rect 33413 33507 33471 33513
rect 33413 33473 33425 33507
rect 33459 33504 33471 33507
rect 33459 33476 34192 33504
rect 33459 33473 33471 33476
rect 33413 33467 33471 33473
rect 27249 33439 27307 33445
rect 27249 33436 27261 33439
rect 26804 33408 27261 33436
rect 26804 33377 26832 33408
rect 27249 33405 27261 33408
rect 27295 33405 27307 33439
rect 27249 33399 27307 33405
rect 27798 33396 27804 33448
rect 27856 33436 27862 33448
rect 28997 33439 29055 33445
rect 28997 33436 29009 33439
rect 27856 33408 29009 33436
rect 27856 33396 27862 33408
rect 28997 33405 29009 33408
rect 29043 33405 29055 33439
rect 28997 33399 29055 33405
rect 33229 33439 33287 33445
rect 33229 33405 33241 33439
rect 33275 33436 33287 33439
rect 34054 33436 34060 33448
rect 33275 33408 34060 33436
rect 33275 33405 33287 33408
rect 33229 33399 33287 33405
rect 34054 33396 34060 33408
rect 34112 33396 34118 33448
rect 34164 33436 34192 33476
rect 34238 33464 34244 33516
rect 34296 33464 34302 33516
rect 34624 33504 34652 33603
rect 36906 33600 36912 33652
rect 36964 33600 36970 33652
rect 34701 33507 34759 33513
rect 34701 33504 34713 33507
rect 34624 33476 34713 33504
rect 34701 33473 34713 33476
rect 34747 33473 34759 33507
rect 34701 33467 34759 33473
rect 36262 33464 36268 33516
rect 36320 33464 36326 33516
rect 36722 33464 36728 33516
rect 36780 33464 36786 33516
rect 36280 33436 36308 33464
rect 34164 33408 36308 33436
rect 26789 33371 26847 33377
rect 26789 33337 26801 33371
rect 26835 33337 26847 33371
rect 26789 33331 26847 33337
rect 33226 33300 33232 33312
rect 26528 33272 33232 33300
rect 33226 33260 33232 33272
rect 33284 33300 33290 33312
rect 34238 33300 34244 33312
rect 33284 33272 34244 33300
rect 33284 33260 33290 33272
rect 34238 33260 34244 33272
rect 34296 33260 34302 33312
rect 34790 33260 34796 33312
rect 34848 33300 34854 33312
rect 34885 33303 34943 33309
rect 34885 33300 34897 33303
rect 34848 33272 34897 33300
rect 34848 33260 34854 33272
rect 34885 33269 34897 33272
rect 34931 33269 34943 33303
rect 34885 33263 34943 33269
rect 1104 33210 38272 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38272 33210
rect 1104 33136 38272 33158
rect 7190 33096 7196 33108
rect 4080 33068 7196 33096
rect 3970 32852 3976 32904
rect 4028 32892 4034 32904
rect 4080 32901 4108 33068
rect 7190 33056 7196 33068
rect 7248 33056 7254 33108
rect 7282 33056 7288 33108
rect 7340 33096 7346 33108
rect 7653 33099 7711 33105
rect 7653 33096 7665 33099
rect 7340 33068 7665 33096
rect 7340 33056 7346 33068
rect 7653 33065 7665 33068
rect 7699 33065 7711 33099
rect 7653 33059 7711 33065
rect 8938 33056 8944 33108
rect 8996 33056 9002 33108
rect 9766 33096 9772 33108
rect 9600 33068 9772 33096
rect 6362 33028 6368 33040
rect 5736 33000 6368 33028
rect 4065 32895 4123 32901
rect 4065 32892 4077 32895
rect 4028 32864 4077 32892
rect 4028 32852 4034 32864
rect 4065 32861 4077 32864
rect 4111 32861 4123 32895
rect 4065 32855 4123 32861
rect 4157 32895 4215 32901
rect 4157 32861 4169 32895
rect 4203 32892 4215 32895
rect 4341 32895 4399 32901
rect 4341 32892 4353 32895
rect 4203 32864 4353 32892
rect 4203 32861 4215 32864
rect 4157 32855 4215 32861
rect 4341 32861 4353 32864
rect 4387 32861 4399 32895
rect 5736 32878 5764 33000
rect 6362 32988 6368 33000
rect 6420 32988 6426 33040
rect 8956 33028 8984 33056
rect 7944 33000 8984 33028
rect 6089 32963 6147 32969
rect 6089 32929 6101 32963
rect 6135 32960 6147 32963
rect 6733 32963 6791 32969
rect 6733 32960 6745 32963
rect 6135 32932 6745 32960
rect 6135 32929 6147 32932
rect 6089 32923 6147 32929
rect 6733 32929 6745 32932
rect 6779 32929 6791 32963
rect 6733 32923 6791 32929
rect 4341 32855 4399 32861
rect 5902 32852 5908 32904
rect 5960 32892 5966 32904
rect 6546 32892 6552 32904
rect 5960 32864 6552 32892
rect 5960 32852 5966 32864
rect 6546 32852 6552 32864
rect 6604 32892 6610 32904
rect 6641 32895 6699 32901
rect 6641 32892 6653 32895
rect 6604 32864 6653 32892
rect 6604 32852 6610 32864
rect 6641 32861 6653 32864
rect 6687 32861 6699 32895
rect 6641 32855 6699 32861
rect 4617 32827 4675 32833
rect 4617 32793 4629 32827
rect 4663 32824 4675 32827
rect 4890 32824 4896 32836
rect 4663 32796 4896 32824
rect 4663 32793 4675 32796
rect 4617 32787 4675 32793
rect 4890 32784 4896 32796
rect 4948 32784 4954 32836
rect 6748 32824 6776 32923
rect 6822 32920 6828 32972
rect 6880 32920 6886 32972
rect 7834 32852 7840 32904
rect 7892 32852 7898 32904
rect 7944 32901 7972 33000
rect 9600 32969 9628 33068
rect 9766 33056 9772 33068
rect 9824 33056 9830 33108
rect 9858 33056 9864 33108
rect 9916 33096 9922 33108
rect 10137 33099 10195 33105
rect 10137 33096 10149 33099
rect 9916 33068 10149 33096
rect 9916 33056 9922 33068
rect 10137 33065 10149 33068
rect 10183 33065 10195 33099
rect 10137 33059 10195 33065
rect 17310 33056 17316 33108
rect 17368 33056 17374 33108
rect 18322 33056 18328 33108
rect 18380 33096 18386 33108
rect 18601 33099 18659 33105
rect 18601 33096 18613 33099
rect 18380 33068 18613 33096
rect 18380 33056 18386 33068
rect 18601 33065 18613 33068
rect 18647 33065 18659 33099
rect 20530 33096 20536 33108
rect 18601 33059 18659 33065
rect 18708 33068 20536 33096
rect 12618 33028 12624 33040
rect 9692 33000 12624 33028
rect 8113 32963 8171 32969
rect 8113 32929 8125 32963
rect 8159 32960 8171 32963
rect 8389 32963 8447 32969
rect 8389 32960 8401 32963
rect 8159 32932 8401 32960
rect 8159 32929 8171 32932
rect 8113 32923 8171 32929
rect 8389 32929 8401 32932
rect 8435 32929 8447 32963
rect 8389 32923 8447 32929
rect 9585 32963 9643 32969
rect 9585 32929 9597 32963
rect 9631 32929 9643 32963
rect 9585 32923 9643 32929
rect 7929 32895 7987 32901
rect 7929 32861 7941 32895
rect 7975 32861 7987 32895
rect 7929 32855 7987 32861
rect 8202 32852 8208 32904
rect 8260 32852 8266 32904
rect 8481 32895 8539 32901
rect 8481 32861 8493 32895
rect 8527 32861 8539 32895
rect 8481 32855 8539 32861
rect 8110 32824 8116 32836
rect 6748 32796 8116 32824
rect 8110 32784 8116 32796
rect 8168 32784 8174 32836
rect 6270 32716 6276 32768
rect 6328 32716 6334 32768
rect 7374 32716 7380 32768
rect 7432 32756 7438 32768
rect 8496 32756 8524 32855
rect 8570 32852 8576 32904
rect 8628 32892 8634 32904
rect 9692 32892 9720 33000
rect 12618 32988 12624 33000
rect 12676 32988 12682 33040
rect 17328 33028 17356 33056
rect 18708 33028 18736 33068
rect 20530 33056 20536 33068
rect 20588 33096 20594 33108
rect 24486 33096 24492 33108
rect 20588 33068 24492 33096
rect 20588 33056 20594 33068
rect 24486 33056 24492 33068
rect 24544 33056 24550 33108
rect 26602 33056 26608 33108
rect 26660 33056 26666 33108
rect 29546 33056 29552 33108
rect 29604 33096 29610 33108
rect 30466 33096 30472 33108
rect 29604 33068 30472 33096
rect 29604 33056 29610 33068
rect 30466 33056 30472 33068
rect 30524 33056 30530 33108
rect 30650 33056 30656 33108
rect 30708 33096 30714 33108
rect 31294 33096 31300 33108
rect 30708 33068 31300 33096
rect 30708 33056 30714 33068
rect 31294 33056 31300 33068
rect 31352 33096 31358 33108
rect 33318 33096 33324 33108
rect 31352 33068 33324 33096
rect 31352 33056 31358 33068
rect 33318 33056 33324 33068
rect 33376 33056 33382 33108
rect 34790 33056 34796 33108
rect 34848 33056 34854 33108
rect 19797 33031 19855 33037
rect 17328 33000 18736 33028
rect 18800 33000 19748 33028
rect 18800 32960 18828 33000
rect 12084 32932 18828 32960
rect 8628 32864 9720 32892
rect 9769 32895 9827 32901
rect 8628 32852 8634 32864
rect 9769 32861 9781 32895
rect 9815 32892 9827 32895
rect 10594 32892 10600 32904
rect 9815 32864 10600 32892
rect 9815 32861 9827 32864
rect 9769 32855 9827 32861
rect 10594 32852 10600 32864
rect 10652 32852 10658 32904
rect 11514 32852 11520 32904
rect 11572 32892 11578 32904
rect 11701 32895 11759 32901
rect 11701 32892 11713 32895
rect 11572 32864 11713 32892
rect 11572 32852 11578 32864
rect 11701 32861 11713 32864
rect 11747 32861 11759 32895
rect 11701 32855 11759 32861
rect 11790 32852 11796 32904
rect 11848 32901 11854 32904
rect 11848 32895 11897 32901
rect 11848 32861 11851 32895
rect 11885 32892 11897 32895
rect 12084 32892 12112 32932
rect 18874 32920 18880 32972
rect 18932 32960 18938 32972
rect 19610 32960 19616 32972
rect 19668 32969 19674 32972
rect 18932 32932 19616 32960
rect 18932 32920 18938 32932
rect 19610 32920 19616 32932
rect 19668 32923 19675 32969
rect 19720 32960 19748 33000
rect 19797 32997 19809 33031
rect 19843 33028 19855 33031
rect 20162 33028 20168 33040
rect 19843 33000 20168 33028
rect 19843 32997 19855 33000
rect 19797 32991 19855 32997
rect 20162 32988 20168 33000
rect 20220 32988 20226 33040
rect 20456 33000 20944 33028
rect 20456 32960 20484 33000
rect 19720 32932 20484 32960
rect 19668 32920 19674 32923
rect 11885 32864 12112 32892
rect 12166 32895 12224 32901
rect 11885 32861 11897 32864
rect 11848 32855 11897 32861
rect 12166 32861 12178 32895
rect 12212 32861 12224 32895
rect 12166 32855 12224 32861
rect 11848 32852 11854 32855
rect 11974 32784 11980 32836
rect 12032 32784 12038 32836
rect 12066 32784 12072 32836
rect 12124 32784 12130 32836
rect 7432 32728 8524 32756
rect 7432 32716 7438 32728
rect 8846 32716 8852 32768
rect 8904 32756 8910 32768
rect 9677 32759 9735 32765
rect 9677 32756 9689 32759
rect 8904 32728 9689 32756
rect 8904 32716 8910 32728
rect 9677 32725 9689 32728
rect 9723 32725 9735 32759
rect 9677 32719 9735 32725
rect 9766 32716 9772 32768
rect 9824 32756 9830 32768
rect 10502 32756 10508 32768
rect 9824 32728 10508 32756
rect 9824 32716 9830 32728
rect 10502 32716 10508 32728
rect 10560 32716 10566 32768
rect 11790 32716 11796 32768
rect 11848 32756 11854 32768
rect 12176 32756 12204 32855
rect 15746 32852 15752 32904
rect 15804 32852 15810 32904
rect 15838 32852 15844 32904
rect 15896 32892 15902 32904
rect 16206 32892 16212 32904
rect 15896 32864 16212 32892
rect 15896 32852 15902 32864
rect 16206 32852 16212 32864
rect 16264 32852 16270 32904
rect 16390 32852 16396 32904
rect 16448 32892 16454 32904
rect 16853 32895 16911 32901
rect 16853 32892 16865 32895
rect 16448 32864 16865 32892
rect 16448 32852 16454 32864
rect 16853 32861 16865 32864
rect 16899 32861 16911 32895
rect 16853 32855 16911 32861
rect 17218 32852 17224 32904
rect 17276 32892 17282 32904
rect 18325 32895 18383 32901
rect 18325 32892 18337 32895
rect 17276 32864 18337 32892
rect 17276 32852 17282 32864
rect 18325 32861 18337 32864
rect 18371 32861 18383 32895
rect 18325 32855 18383 32861
rect 18690 32852 18696 32904
rect 18748 32852 18754 32904
rect 19702 32892 19708 32904
rect 19628 32864 19708 32892
rect 15764 32824 15792 32852
rect 18230 32824 18236 32836
rect 15764 32796 18236 32824
rect 18230 32784 18236 32796
rect 18288 32824 18294 32836
rect 18417 32827 18475 32833
rect 18417 32824 18429 32827
rect 18288 32796 18429 32824
rect 18288 32784 18294 32796
rect 18417 32793 18429 32796
rect 18463 32793 18475 32827
rect 18417 32787 18475 32793
rect 18785 32827 18843 32833
rect 18785 32793 18797 32827
rect 18831 32824 18843 32827
rect 19058 32824 19064 32836
rect 18831 32796 19064 32824
rect 18831 32793 18843 32796
rect 18785 32787 18843 32793
rect 11848 32728 12204 32756
rect 11848 32716 11854 32728
rect 12342 32716 12348 32768
rect 12400 32716 12406 32768
rect 16393 32759 16451 32765
rect 16393 32725 16405 32759
rect 16439 32756 16451 32759
rect 16666 32756 16672 32768
rect 16439 32728 16672 32756
rect 16439 32725 16451 32728
rect 16393 32719 16451 32725
rect 16666 32716 16672 32728
rect 16724 32716 16730 32768
rect 18432 32756 18460 32787
rect 19058 32784 19064 32796
rect 19116 32784 19122 32836
rect 19628 32833 19656 32864
rect 19702 32852 19708 32864
rect 19760 32852 19766 32904
rect 19889 32895 19947 32901
rect 19889 32861 19901 32895
rect 19935 32861 19947 32895
rect 19889 32855 19947 32861
rect 20165 32895 20223 32901
rect 20165 32861 20177 32895
rect 20211 32892 20223 32895
rect 20254 32892 20260 32904
rect 20211 32864 20260 32892
rect 20211 32861 20223 32864
rect 20165 32855 20223 32861
rect 19613 32827 19671 32833
rect 19613 32793 19625 32827
rect 19659 32793 19671 32827
rect 19613 32787 19671 32793
rect 19904 32756 19932 32855
rect 20254 32852 20260 32864
rect 20312 32852 20318 32904
rect 20456 32901 20484 32932
rect 20916 32904 20944 33000
rect 22002 32988 22008 33040
rect 22060 33028 22066 33040
rect 26142 33028 26148 33040
rect 22060 33000 26148 33028
rect 22060 32988 22066 33000
rect 22020 32960 22048 32988
rect 22296 32969 22324 33000
rect 26142 32988 26148 33000
rect 26200 32988 26206 33040
rect 21836 32932 22048 32960
rect 22281 32963 22339 32969
rect 20441 32895 20499 32901
rect 20441 32861 20453 32895
rect 20487 32861 20499 32895
rect 20441 32855 20499 32861
rect 20530 32852 20536 32904
rect 20588 32852 20594 32904
rect 20898 32852 20904 32904
rect 20956 32852 20962 32904
rect 21450 32852 21456 32904
rect 21508 32852 21514 32904
rect 19978 32784 19984 32836
rect 20036 32824 20042 32836
rect 20349 32827 20407 32833
rect 20349 32824 20361 32827
rect 20036 32796 20361 32824
rect 20036 32784 20042 32796
rect 20349 32793 20361 32796
rect 20395 32824 20407 32827
rect 21836 32824 21864 32932
rect 22281 32929 22293 32963
rect 22327 32929 22339 32963
rect 22281 32923 22339 32929
rect 26878 32920 26884 32972
rect 26936 32960 26942 32972
rect 27157 32963 27215 32969
rect 27157 32960 27169 32963
rect 26936 32932 27169 32960
rect 26936 32920 26942 32932
rect 27157 32929 27169 32932
rect 27203 32929 27215 32963
rect 27798 32960 27804 32972
rect 27157 32923 27215 32929
rect 27448 32932 27804 32960
rect 21910 32852 21916 32904
rect 21968 32892 21974 32904
rect 22097 32895 22155 32901
rect 22097 32892 22109 32895
rect 21968 32864 22109 32892
rect 21968 32852 21974 32864
rect 22097 32861 22109 32864
rect 22143 32892 22155 32895
rect 22186 32892 22192 32904
rect 22143 32864 22192 32892
rect 22143 32861 22155 32864
rect 22097 32855 22155 32861
rect 22186 32852 22192 32864
rect 22244 32852 22250 32904
rect 22830 32852 22836 32904
rect 22888 32892 22894 32904
rect 23385 32895 23443 32901
rect 23385 32892 23397 32895
rect 22888 32864 23397 32892
rect 22888 32852 22894 32864
rect 23385 32861 23397 32864
rect 23431 32861 23443 32895
rect 27448 32892 27476 32932
rect 27798 32920 27804 32932
rect 27856 32920 27862 32972
rect 28534 32920 28540 32972
rect 28592 32960 28598 32972
rect 34808 32960 34836 33056
rect 34977 32963 35035 32969
rect 34977 32960 34989 32963
rect 28592 32932 28856 32960
rect 28592 32920 28598 32932
rect 28828 32904 28856 32932
rect 30392 32932 33548 32960
rect 34808 32932 34989 32960
rect 23385 32855 23443 32861
rect 26988 32864 27476 32892
rect 23201 32827 23259 32833
rect 23201 32824 23213 32827
rect 20395 32796 21864 32824
rect 22388 32796 23213 32824
rect 20395 32793 20407 32796
rect 20349 32787 20407 32793
rect 18432 32728 19932 32756
rect 20714 32716 20720 32768
rect 20772 32716 20778 32768
rect 21542 32716 21548 32768
rect 21600 32756 21606 32768
rect 22388 32756 22416 32796
rect 23201 32793 23213 32796
rect 23247 32793 23259 32827
rect 23201 32787 23259 32793
rect 21600 32728 22416 32756
rect 23569 32759 23627 32765
rect 21600 32716 21606 32728
rect 23569 32725 23581 32759
rect 23615 32756 23627 32759
rect 23934 32756 23940 32768
rect 23615 32728 23940 32756
rect 23615 32725 23627 32728
rect 23569 32719 23627 32725
rect 23934 32716 23940 32728
rect 23992 32716 23998 32768
rect 26326 32716 26332 32768
rect 26384 32756 26390 32768
rect 26602 32756 26608 32768
rect 26384 32728 26608 32756
rect 26384 32716 26390 32728
rect 26602 32716 26608 32728
rect 26660 32756 26666 32768
rect 26988 32765 27016 32864
rect 27522 32852 27528 32904
rect 27580 32852 27586 32904
rect 28810 32852 28816 32904
rect 28868 32892 28874 32904
rect 30282 32892 30288 32904
rect 28868 32864 28934 32892
rect 29104 32864 30288 32892
rect 28868 32852 28874 32864
rect 29104 32836 29132 32864
rect 30282 32852 30288 32864
rect 30340 32892 30346 32904
rect 30392 32901 30420 32932
rect 30377 32895 30435 32901
rect 30377 32892 30389 32895
rect 30340 32864 30389 32892
rect 30340 32852 30346 32864
rect 30377 32861 30389 32864
rect 30423 32861 30435 32895
rect 30377 32855 30435 32861
rect 30926 32852 30932 32904
rect 30984 32852 30990 32904
rect 31202 32852 31208 32904
rect 31260 32852 31266 32904
rect 32490 32852 32496 32904
rect 32548 32892 32554 32904
rect 32950 32892 32956 32904
rect 32548 32864 32956 32892
rect 32548 32852 32554 32864
rect 32950 32852 32956 32864
rect 33008 32852 33014 32904
rect 33520 32892 33548 32932
rect 34977 32929 34989 32932
rect 35023 32929 35035 32963
rect 34977 32923 35035 32929
rect 34330 32892 34336 32904
rect 33520 32864 34336 32892
rect 34330 32852 34336 32864
rect 34388 32852 34394 32904
rect 34425 32895 34483 32901
rect 34425 32861 34437 32895
rect 34471 32892 34483 32895
rect 34701 32895 34759 32901
rect 34701 32892 34713 32895
rect 34471 32864 34713 32892
rect 34471 32861 34483 32864
rect 34425 32855 34483 32861
rect 34701 32861 34713 32864
rect 34747 32861 34759 32895
rect 34701 32855 34759 32861
rect 35986 32852 35992 32904
rect 36044 32892 36050 32904
rect 36044 32864 36110 32892
rect 36044 32852 36050 32864
rect 27801 32827 27859 32833
rect 27801 32793 27813 32827
rect 27847 32824 27859 32827
rect 28074 32824 28080 32836
rect 27847 32796 28080 32824
rect 27847 32793 27859 32796
rect 27801 32787 27859 32793
rect 28074 32784 28080 32796
rect 28132 32784 28138 32836
rect 29086 32784 29092 32836
rect 29144 32784 29150 32836
rect 31481 32827 31539 32833
rect 31481 32793 31493 32827
rect 31527 32793 31539 32827
rect 31481 32787 31539 32793
rect 36725 32827 36783 32833
rect 36725 32793 36737 32827
rect 36771 32793 36783 32827
rect 36725 32787 36783 32793
rect 26973 32759 27031 32765
rect 26973 32756 26985 32759
rect 26660 32728 26985 32756
rect 26660 32716 26666 32728
rect 26973 32725 26985 32728
rect 27019 32725 27031 32759
rect 26973 32719 27031 32725
rect 27065 32759 27123 32765
rect 27065 32725 27077 32759
rect 27111 32756 27123 32759
rect 27246 32756 27252 32768
rect 27111 32728 27252 32756
rect 27111 32725 27123 32728
rect 27065 32719 27123 32725
rect 27246 32716 27252 32728
rect 27304 32756 27310 32768
rect 27614 32756 27620 32768
rect 27304 32728 27620 32756
rect 27304 32716 27310 32728
rect 27614 32716 27620 32728
rect 27672 32716 27678 32768
rect 28718 32716 28724 32768
rect 28776 32756 28782 32768
rect 29273 32759 29331 32765
rect 29273 32756 29285 32759
rect 28776 32728 29285 32756
rect 28776 32716 28782 32728
rect 29273 32725 29285 32728
rect 29319 32725 29331 32759
rect 29273 32719 29331 32725
rect 30190 32716 30196 32768
rect 30248 32716 30254 32768
rect 31113 32759 31171 32765
rect 31113 32725 31125 32759
rect 31159 32756 31171 32759
rect 31496 32756 31524 32787
rect 31159 32728 31524 32756
rect 31159 32725 31171 32728
rect 31113 32719 31171 32725
rect 32122 32716 32128 32768
rect 32180 32756 32186 32768
rect 32953 32759 33011 32765
rect 32953 32756 32965 32759
rect 32180 32728 32965 32756
rect 32180 32716 32186 32728
rect 32953 32725 32965 32728
rect 32999 32725 33011 32759
rect 32953 32719 33011 32725
rect 35618 32716 35624 32768
rect 35676 32756 35682 32768
rect 36740 32756 36768 32787
rect 35676 32728 36768 32756
rect 35676 32716 35682 32728
rect 1104 32666 38272 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38272 32666
rect 1104 32592 38272 32614
rect 4890 32512 4896 32564
rect 4948 32552 4954 32564
rect 4985 32555 5043 32561
rect 4985 32552 4997 32555
rect 4948 32524 4997 32552
rect 4948 32512 4954 32524
rect 4985 32521 4997 32524
rect 5031 32521 5043 32555
rect 4985 32515 5043 32521
rect 6270 32512 6276 32564
rect 6328 32512 6334 32564
rect 8110 32512 8116 32564
rect 8168 32512 8174 32564
rect 12069 32555 12127 32561
rect 12069 32521 12081 32555
rect 12115 32521 12127 32555
rect 12069 32515 12127 32521
rect 5169 32419 5227 32425
rect 5169 32385 5181 32419
rect 5215 32416 5227 32419
rect 6288 32416 6316 32512
rect 8128 32484 8156 32512
rect 11793 32487 11851 32493
rect 11793 32484 11805 32487
rect 8128 32456 11805 32484
rect 11793 32453 11805 32456
rect 11839 32484 11851 32487
rect 12084 32484 12112 32515
rect 12342 32512 12348 32564
rect 12400 32552 12406 32564
rect 16853 32555 16911 32561
rect 16853 32552 16865 32555
rect 12400 32524 12480 32552
rect 12400 32512 12406 32524
rect 12452 32493 12480 32524
rect 16408 32524 16865 32552
rect 16408 32496 16436 32524
rect 16853 32521 16865 32524
rect 16899 32521 16911 32555
rect 16853 32515 16911 32521
rect 17678 32512 17684 32564
rect 17736 32512 17742 32564
rect 23382 32552 23388 32564
rect 17880 32524 22232 32552
rect 12253 32487 12311 32493
rect 12253 32484 12265 32487
rect 11839 32456 12020 32484
rect 12084 32456 12265 32484
rect 11839 32453 11851 32456
rect 11793 32447 11851 32453
rect 5215 32388 6316 32416
rect 11517 32419 11575 32425
rect 5215 32385 5227 32388
rect 5169 32379 5227 32385
rect 11517 32385 11529 32419
rect 11563 32416 11575 32419
rect 11701 32419 11759 32425
rect 11563 32388 11652 32416
rect 11563 32385 11575 32388
rect 11517 32379 11575 32385
rect 5718 32308 5724 32360
rect 5776 32348 5782 32360
rect 8294 32348 8300 32360
rect 5776 32320 8300 32348
rect 5776 32308 5782 32320
rect 8294 32308 8300 32320
rect 8352 32308 8358 32360
rect 11624 32224 11652 32388
rect 11701 32385 11713 32419
rect 11747 32385 11759 32419
rect 11701 32379 11759 32385
rect 11716 32280 11744 32379
rect 11882 32376 11888 32428
rect 11940 32376 11946 32428
rect 11992 32416 12020 32456
rect 12253 32453 12265 32456
rect 12299 32453 12311 32487
rect 12253 32447 12311 32453
rect 12437 32487 12495 32493
rect 12437 32453 12449 32487
rect 12483 32453 12495 32487
rect 12437 32447 12495 32453
rect 16390 32444 16396 32496
rect 16448 32444 16454 32496
rect 16669 32487 16727 32493
rect 16669 32453 16681 32487
rect 16715 32484 16727 32487
rect 17034 32484 17040 32496
rect 16715 32456 17040 32484
rect 16715 32453 16727 32456
rect 16669 32447 16727 32453
rect 17034 32444 17040 32456
rect 17092 32484 17098 32496
rect 17313 32487 17371 32493
rect 17313 32484 17325 32487
rect 17092 32456 17325 32484
rect 17092 32444 17098 32456
rect 17313 32453 17325 32456
rect 17359 32453 17371 32487
rect 17313 32447 17371 32453
rect 17494 32444 17500 32496
rect 17552 32444 17558 32496
rect 13538 32416 13544 32428
rect 11992 32388 13544 32416
rect 13538 32376 13544 32388
rect 13596 32376 13602 32428
rect 17880 32416 17908 32524
rect 20254 32444 20260 32496
rect 20312 32484 20318 32496
rect 21634 32484 21640 32496
rect 20312 32456 21640 32484
rect 20312 32444 20318 32456
rect 21634 32444 21640 32456
rect 21692 32444 21698 32496
rect 17512 32388 17908 32416
rect 16114 32308 16120 32360
rect 16172 32308 16178 32360
rect 12250 32280 12256 32292
rect 11716 32252 12256 32280
rect 12250 32240 12256 32252
rect 12308 32240 12314 32292
rect 12621 32283 12679 32289
rect 12621 32249 12633 32283
rect 12667 32280 12679 32283
rect 13630 32280 13636 32292
rect 12667 32252 13636 32280
rect 12667 32249 12679 32252
rect 12621 32243 12679 32249
rect 13630 32240 13636 32252
rect 13688 32240 13694 32292
rect 16132 32280 16160 32308
rect 17037 32283 17095 32289
rect 17037 32280 17049 32283
rect 16132 32252 17049 32280
rect 17037 32249 17049 32252
rect 17083 32280 17095 32283
rect 17512 32280 17540 32388
rect 18414 32376 18420 32428
rect 18472 32376 18478 32428
rect 18598 32376 18604 32428
rect 18656 32376 18662 32428
rect 18690 32376 18696 32428
rect 18748 32376 18754 32428
rect 18877 32419 18935 32425
rect 18877 32385 18889 32419
rect 18923 32385 18935 32419
rect 18877 32379 18935 32385
rect 18892 32348 18920 32379
rect 18966 32376 18972 32428
rect 19024 32376 19030 32428
rect 19058 32376 19064 32428
rect 19116 32376 19122 32428
rect 19076 32348 19104 32376
rect 18892 32320 19104 32348
rect 17083 32252 17540 32280
rect 17083 32249 17095 32252
rect 17037 32243 17095 32249
rect 17586 32240 17592 32292
rect 17644 32280 17650 32292
rect 20272 32280 20300 32444
rect 21266 32376 21272 32428
rect 21324 32376 21330 32428
rect 21358 32376 21364 32428
rect 21416 32416 21422 32428
rect 21913 32419 21971 32425
rect 21913 32416 21925 32419
rect 21416 32388 21925 32416
rect 21416 32376 21422 32388
rect 21913 32385 21925 32388
rect 21959 32385 21971 32419
rect 21913 32379 21971 32385
rect 17644 32252 20300 32280
rect 22204 32280 22232 32524
rect 22756 32524 23388 32552
rect 22278 32376 22284 32428
rect 22336 32416 22342 32428
rect 22756 32416 22784 32524
rect 23382 32512 23388 32524
rect 23440 32512 23446 32564
rect 23842 32512 23848 32564
rect 23900 32552 23906 32564
rect 23900 32524 26004 32552
rect 23900 32512 23906 32524
rect 22830 32444 22836 32496
rect 22888 32484 22894 32496
rect 23109 32487 23167 32493
rect 23109 32484 23121 32487
rect 22888 32456 23121 32484
rect 22888 32444 22894 32456
rect 23109 32453 23121 32456
rect 23155 32453 23167 32487
rect 23109 32447 23167 32453
rect 23201 32487 23259 32493
rect 23201 32453 23213 32487
rect 23247 32484 23259 32487
rect 23290 32484 23296 32496
rect 23247 32456 23296 32484
rect 23247 32453 23259 32456
rect 23201 32447 23259 32453
rect 23290 32444 23296 32456
rect 23348 32444 23354 32496
rect 23017 32419 23075 32425
rect 23017 32416 23029 32419
rect 22336 32388 23029 32416
rect 22336 32376 22342 32388
rect 23017 32385 23029 32388
rect 23063 32385 23075 32419
rect 23017 32379 23075 32385
rect 23382 32376 23388 32428
rect 23440 32376 23446 32428
rect 23753 32419 23811 32425
rect 23753 32385 23765 32419
rect 23799 32416 23811 32419
rect 23860 32416 23888 32512
rect 23934 32444 23940 32496
rect 23992 32444 23998 32496
rect 25976 32428 26004 32524
rect 27522 32512 27528 32564
rect 27580 32552 27586 32564
rect 27801 32555 27859 32561
rect 27801 32552 27813 32555
rect 27580 32524 27813 32552
rect 27580 32512 27586 32524
rect 27801 32521 27813 32524
rect 27847 32521 27859 32555
rect 27801 32515 27859 32521
rect 28074 32512 28080 32564
rect 28132 32552 28138 32564
rect 28997 32555 29055 32561
rect 28997 32552 29009 32555
rect 28132 32524 29009 32552
rect 28132 32512 28138 32524
rect 28997 32521 29009 32524
rect 29043 32521 29055 32555
rect 28997 32515 29055 32521
rect 31202 32512 31208 32564
rect 31260 32552 31266 32564
rect 31389 32555 31447 32561
rect 31389 32552 31401 32555
rect 31260 32524 31401 32552
rect 31260 32512 31266 32524
rect 31389 32521 31401 32524
rect 31435 32521 31447 32555
rect 31389 32515 31447 32521
rect 35989 32555 36047 32561
rect 35989 32521 36001 32555
rect 36035 32552 36047 32555
rect 36722 32552 36728 32564
rect 36035 32524 36728 32552
rect 36035 32521 36047 32524
rect 35989 32515 36047 32521
rect 36722 32512 36728 32524
rect 36780 32512 36786 32564
rect 27706 32444 27712 32496
rect 27764 32484 27770 32496
rect 32582 32484 32588 32496
rect 27764 32456 32588 32484
rect 27764 32444 27770 32456
rect 23799 32388 23888 32416
rect 24029 32419 24087 32425
rect 23799 32385 23811 32388
rect 23753 32379 23811 32385
rect 24029 32385 24041 32419
rect 24075 32385 24087 32419
rect 24029 32379 24087 32385
rect 23106 32308 23112 32360
rect 23164 32348 23170 32360
rect 24044 32348 24072 32379
rect 24118 32376 24124 32428
rect 24176 32376 24182 32428
rect 25958 32376 25964 32428
rect 26016 32376 26022 32428
rect 27724 32416 27752 32444
rect 27893 32419 27951 32425
rect 27893 32416 27905 32419
rect 27724 32388 27905 32416
rect 27893 32385 27905 32388
rect 27939 32385 27951 32419
rect 27893 32379 27951 32385
rect 28537 32419 28595 32425
rect 28537 32385 28549 32419
rect 28583 32416 28595 32419
rect 28718 32416 28724 32428
rect 28583 32388 28724 32416
rect 28583 32385 28595 32388
rect 28537 32379 28595 32385
rect 23164 32320 24072 32348
rect 23164 32308 23170 32320
rect 24762 32308 24768 32360
rect 24820 32308 24826 32360
rect 25774 32308 25780 32360
rect 25832 32348 25838 32360
rect 25832 32320 26464 32348
rect 25832 32308 25838 32320
rect 24780 32280 24808 32308
rect 22204 32252 24808 32280
rect 17644 32240 17650 32252
rect 11606 32172 11612 32224
rect 11664 32172 11670 32224
rect 15654 32172 15660 32224
rect 15712 32212 15718 32224
rect 16758 32212 16764 32224
rect 15712 32184 16764 32212
rect 15712 32172 15718 32184
rect 16758 32172 16764 32184
rect 16816 32212 16822 32224
rect 16853 32215 16911 32221
rect 16853 32212 16865 32215
rect 16816 32184 16865 32212
rect 16816 32172 16822 32184
rect 16853 32181 16865 32184
rect 16899 32212 16911 32215
rect 17126 32212 17132 32224
rect 16899 32184 17132 32212
rect 16899 32181 16911 32184
rect 16853 32175 16911 32181
rect 17126 32172 17132 32184
rect 17184 32212 17190 32224
rect 17497 32215 17555 32221
rect 17497 32212 17509 32215
rect 17184 32184 17509 32212
rect 17184 32172 17190 32184
rect 17497 32181 17509 32184
rect 17543 32212 17555 32215
rect 19426 32212 19432 32224
rect 17543 32184 19432 32212
rect 17543 32181 17555 32184
rect 17497 32175 17555 32181
rect 19426 32172 19432 32184
rect 19484 32172 19490 32224
rect 19978 32172 19984 32224
rect 20036 32172 20042 32224
rect 22186 32172 22192 32224
rect 22244 32172 22250 32224
rect 22830 32172 22836 32224
rect 22888 32172 22894 32224
rect 24305 32215 24363 32221
rect 24305 32181 24317 32215
rect 24351 32212 24363 32215
rect 25314 32212 25320 32224
rect 24351 32184 25320 32212
rect 24351 32181 24363 32184
rect 24305 32175 24363 32181
rect 25314 32172 25320 32184
rect 25372 32172 25378 32224
rect 26436 32212 26464 32320
rect 27982 32308 27988 32360
rect 28040 32348 28046 32360
rect 28261 32351 28319 32357
rect 28261 32348 28273 32351
rect 28040 32320 28273 32348
rect 28040 32308 28046 32320
rect 28261 32317 28273 32320
rect 28307 32348 28319 32351
rect 28350 32348 28356 32360
rect 28307 32320 28356 32348
rect 28307 32317 28319 32320
rect 28261 32311 28319 32317
rect 28350 32308 28356 32320
rect 28408 32308 28414 32360
rect 28442 32308 28448 32360
rect 28500 32308 28506 32360
rect 26694 32240 26700 32292
rect 26752 32280 26758 32292
rect 28552 32280 28580 32379
rect 28718 32376 28724 32388
rect 28776 32376 28782 32428
rect 29181 32419 29239 32425
rect 29181 32416 29193 32419
rect 28920 32388 29193 32416
rect 28920 32289 28948 32388
rect 29181 32385 29193 32388
rect 29227 32385 29239 32419
rect 29181 32379 29239 32385
rect 30745 32419 30803 32425
rect 30745 32385 30757 32419
rect 30791 32385 30803 32419
rect 30745 32379 30803 32385
rect 30650 32308 30656 32360
rect 30708 32308 30714 32360
rect 30760 32348 30788 32379
rect 30834 32376 30840 32428
rect 30892 32376 30898 32428
rect 31496 32425 31524 32456
rect 32582 32444 32588 32456
rect 32640 32484 32646 32496
rect 34606 32484 34612 32496
rect 32640 32456 34612 32484
rect 32640 32444 32646 32456
rect 34606 32444 34612 32456
rect 34664 32444 34670 32496
rect 31481 32419 31539 32425
rect 31481 32385 31493 32419
rect 31527 32385 31539 32419
rect 32122 32416 32128 32428
rect 31481 32379 31539 32385
rect 31726 32388 32128 32416
rect 31726 32348 31754 32388
rect 32122 32376 32128 32388
rect 32180 32376 32186 32428
rect 32214 32376 32220 32428
rect 32272 32416 32278 32428
rect 32401 32419 32459 32425
rect 32401 32416 32413 32419
rect 32272 32388 32413 32416
rect 32272 32376 32278 32388
rect 32401 32385 32413 32388
rect 32447 32385 32459 32419
rect 32401 32379 32459 32385
rect 33134 32376 33140 32428
rect 33192 32376 33198 32428
rect 33226 32376 33232 32428
rect 33284 32416 33290 32428
rect 33413 32419 33471 32425
rect 33413 32416 33425 32419
rect 33284 32388 33425 32416
rect 33284 32376 33290 32388
rect 33413 32385 33425 32388
rect 33459 32416 33471 32419
rect 35618 32416 35624 32428
rect 33459 32388 35624 32416
rect 33459 32385 33471 32388
rect 33413 32379 33471 32385
rect 35618 32376 35624 32388
rect 35676 32376 35682 32428
rect 35805 32419 35863 32425
rect 35805 32385 35817 32419
rect 35851 32385 35863 32419
rect 35805 32379 35863 32385
rect 30760 32320 31754 32348
rect 32306 32308 32312 32360
rect 32364 32348 32370 32360
rect 32677 32351 32735 32357
rect 32677 32348 32689 32351
rect 32364 32320 32689 32348
rect 32364 32308 32370 32320
rect 32677 32317 32689 32320
rect 32723 32317 32735 32351
rect 32677 32311 32735 32317
rect 26752 32252 28580 32280
rect 28905 32283 28963 32289
rect 26752 32240 26758 32252
rect 28905 32249 28917 32283
rect 28951 32249 28963 32283
rect 28905 32243 28963 32249
rect 30926 32240 30932 32292
rect 30984 32280 30990 32292
rect 31205 32283 31263 32289
rect 31205 32280 31217 32283
rect 30984 32252 31217 32280
rect 30984 32240 30990 32252
rect 31205 32249 31217 32252
rect 31251 32249 31263 32283
rect 31205 32243 31263 32249
rect 32858 32240 32864 32292
rect 32916 32240 32922 32292
rect 35820 32212 35848 32379
rect 26436 32184 35848 32212
rect 1104 32122 38272 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38272 32122
rect 1104 32048 38272 32070
rect 4512 32011 4570 32017
rect 4512 31977 4524 32011
rect 4558 32008 4570 32011
rect 7285 32011 7343 32017
rect 7285 32008 7297 32011
rect 4558 31980 7297 32008
rect 4558 31977 4570 31980
rect 4512 31971 4570 31977
rect 7285 31977 7297 31980
rect 7331 31977 7343 32011
rect 7285 31971 7343 31977
rect 7834 31968 7840 32020
rect 7892 32008 7898 32020
rect 8570 32008 8576 32020
rect 7892 31980 8576 32008
rect 7892 31968 7898 31980
rect 8570 31968 8576 31980
rect 8628 31968 8634 32020
rect 9600 31980 11652 32008
rect 9600 31940 9628 31980
rect 11624 31952 11652 31980
rect 13538 31968 13544 32020
rect 13596 32008 13602 32020
rect 17586 32008 17592 32020
rect 13596 31980 17592 32008
rect 13596 31968 13602 31980
rect 17586 31968 17592 31980
rect 17644 31968 17650 32020
rect 18138 31968 18144 32020
rect 18196 32008 18202 32020
rect 18966 32008 18972 32020
rect 18196 31980 18972 32008
rect 18196 31968 18202 31980
rect 18966 31968 18972 31980
rect 19024 31968 19030 32020
rect 19058 31968 19064 32020
rect 19116 31968 19122 32020
rect 22002 31968 22008 32020
rect 22060 32008 22066 32020
rect 22554 32008 22560 32020
rect 22060 31980 22560 32008
rect 22060 31968 22066 31980
rect 22554 31968 22560 31980
rect 22612 31968 22618 32020
rect 24029 32011 24087 32017
rect 22664 31980 23152 32008
rect 6656 31912 9628 31940
rect 5718 31832 5724 31884
rect 5776 31832 5782 31884
rect 6656 31881 6684 31912
rect 11606 31900 11612 31952
rect 11664 31940 11670 31952
rect 11664 31912 19334 31940
rect 11664 31900 11670 31912
rect 6273 31875 6331 31881
rect 6273 31841 6285 31875
rect 6319 31872 6331 31875
rect 6641 31875 6699 31881
rect 6641 31872 6653 31875
rect 6319 31844 6653 31872
rect 6319 31841 6331 31844
rect 6273 31835 6331 31841
rect 6641 31841 6653 31844
rect 6687 31841 6699 31875
rect 6641 31835 6699 31841
rect 7193 31875 7251 31881
rect 7193 31841 7205 31875
rect 7239 31872 7251 31875
rect 7239 31844 7880 31872
rect 7239 31841 7251 31844
rect 7193 31835 7251 31841
rect 3970 31764 3976 31816
rect 4028 31764 4034 31816
rect 4065 31807 4123 31813
rect 4065 31773 4077 31807
rect 4111 31804 4123 31807
rect 4249 31807 4307 31813
rect 4249 31804 4261 31807
rect 4111 31776 4261 31804
rect 4111 31773 4123 31776
rect 4065 31767 4123 31773
rect 4249 31773 4261 31776
rect 4295 31773 4307 31807
rect 5736 31804 5764 31832
rect 5658 31776 5764 31804
rect 4249 31767 4307 31773
rect 6546 31764 6552 31816
rect 6604 31804 6610 31816
rect 6604 31776 7052 31804
rect 6604 31764 6610 31776
rect 7024 31736 7052 31776
rect 7374 31764 7380 31816
rect 7432 31804 7438 31816
rect 7469 31807 7527 31813
rect 7469 31804 7481 31807
rect 7432 31776 7481 31804
rect 7432 31764 7438 31776
rect 7469 31773 7481 31776
rect 7515 31773 7527 31807
rect 7469 31767 7527 31773
rect 7561 31807 7619 31813
rect 7561 31773 7573 31807
rect 7607 31773 7619 31807
rect 7561 31767 7619 31773
rect 7576 31736 7604 31767
rect 7650 31764 7656 31816
rect 7708 31764 7714 31816
rect 7852 31813 7880 31844
rect 8036 31844 8892 31872
rect 7837 31807 7895 31813
rect 7837 31773 7849 31807
rect 7883 31773 7895 31807
rect 8036 31804 8064 31844
rect 8864 31816 8892 31844
rect 9030 31832 9036 31884
rect 9088 31872 9094 31884
rect 9088 31844 9260 31872
rect 9088 31832 9094 31844
rect 7837 31767 7895 31773
rect 7944 31776 8064 31804
rect 7944 31736 7972 31776
rect 8110 31764 8116 31816
rect 8168 31764 8174 31816
rect 8478 31764 8484 31816
rect 8536 31764 8542 31816
rect 8846 31764 8852 31816
rect 8904 31764 8910 31816
rect 9232 31813 9260 31844
rect 17954 31832 17960 31884
rect 18012 31832 18018 31884
rect 18322 31832 18328 31884
rect 18380 31872 18386 31884
rect 19306 31872 19334 31912
rect 20346 31900 20352 31952
rect 20404 31940 20410 31952
rect 21818 31940 21824 31952
rect 20404 31912 21824 31940
rect 20404 31900 20410 31912
rect 21818 31900 21824 31912
rect 21876 31900 21882 31952
rect 20622 31872 20628 31884
rect 18380 31844 19104 31872
rect 19306 31844 20628 31872
rect 18380 31832 18386 31844
rect 9217 31807 9275 31813
rect 9217 31773 9229 31807
rect 9263 31773 9275 31807
rect 9217 31767 9275 31773
rect 9309 31807 9367 31813
rect 9309 31773 9321 31807
rect 9355 31804 9367 31807
rect 9493 31807 9551 31813
rect 9493 31804 9505 31807
rect 9355 31776 9505 31804
rect 9355 31773 9367 31776
rect 9309 31767 9367 31773
rect 9493 31773 9505 31776
rect 9539 31773 9551 31807
rect 9493 31767 9551 31773
rect 13633 31807 13691 31813
rect 13633 31773 13645 31807
rect 13679 31804 13691 31807
rect 14458 31804 14464 31816
rect 13679 31776 14464 31804
rect 13679 31773 13691 31776
rect 13633 31767 13691 31773
rect 14458 31764 14464 31776
rect 14516 31764 14522 31816
rect 15470 31764 15476 31816
rect 15528 31804 15534 31816
rect 16390 31804 16396 31816
rect 15528 31776 16396 31804
rect 15528 31764 15534 31776
rect 16390 31764 16396 31776
rect 16448 31804 16454 31816
rect 17972 31804 18000 31832
rect 19076 31813 19104 31844
rect 20622 31832 20628 31844
rect 20680 31872 20686 31884
rect 22664 31872 22692 31980
rect 23124 31952 23152 31980
rect 24029 31977 24041 32011
rect 24075 32008 24087 32011
rect 24075 31980 25084 32008
rect 24075 31977 24087 31980
rect 24029 31971 24087 31977
rect 22738 31900 22744 31952
rect 22796 31940 22802 31952
rect 23014 31940 23020 31952
rect 22796 31912 23020 31940
rect 22796 31900 22802 31912
rect 23014 31900 23020 31912
rect 23072 31900 23078 31952
rect 23106 31900 23112 31952
rect 23164 31900 23170 31952
rect 23382 31900 23388 31952
rect 23440 31940 23446 31952
rect 24949 31943 25007 31949
rect 23440 31912 24532 31940
rect 23440 31900 23446 31912
rect 24118 31872 24124 31884
rect 20680 31844 22692 31872
rect 22996 31844 23520 31872
rect 20680 31832 20686 31844
rect 18877 31807 18935 31813
rect 18877 31804 18889 31807
rect 16448 31776 16712 31804
rect 17972 31776 18889 31804
rect 16448 31764 16454 31776
rect 7024 31708 7972 31736
rect 9766 31696 9772 31748
rect 9824 31696 9830 31748
rect 10318 31696 10324 31748
rect 10376 31696 10382 31748
rect 12894 31696 12900 31748
rect 12952 31736 12958 31748
rect 13081 31739 13139 31745
rect 13081 31736 13093 31739
rect 12952 31708 13093 31736
rect 12952 31696 12958 31708
rect 13081 31705 13093 31708
rect 13127 31705 13139 31739
rect 13081 31699 13139 31705
rect 13262 31696 13268 31748
rect 13320 31696 13326 31748
rect 13906 31736 13912 31748
rect 13464 31708 13912 31736
rect 7834 31628 7840 31680
rect 7892 31668 7898 31680
rect 8021 31671 8079 31677
rect 8021 31668 8033 31671
rect 7892 31640 8033 31668
rect 7892 31628 7898 31640
rect 8021 31637 8033 31640
rect 8067 31637 8079 31671
rect 8021 31631 8079 31637
rect 8294 31628 8300 31680
rect 8352 31628 8358 31680
rect 11241 31671 11299 31677
rect 11241 31637 11253 31671
rect 11287 31668 11299 31671
rect 11606 31668 11612 31680
rect 11287 31640 11612 31668
rect 11287 31637 11299 31640
rect 11241 31631 11299 31637
rect 11606 31628 11612 31640
rect 11664 31628 11670 31680
rect 13354 31628 13360 31680
rect 13412 31628 13418 31680
rect 13464 31677 13492 31708
rect 13906 31696 13912 31708
rect 13964 31696 13970 31748
rect 13449 31671 13507 31677
rect 13449 31637 13461 31671
rect 13495 31637 13507 31671
rect 16684 31668 16712 31776
rect 18877 31773 18889 31776
rect 18923 31773 18935 31807
rect 18877 31767 18935 31773
rect 19061 31807 19119 31813
rect 19061 31773 19073 31807
rect 19107 31773 19119 31807
rect 19061 31767 19119 31773
rect 21266 31764 21272 31816
rect 21324 31764 21330 31816
rect 21910 31764 21916 31816
rect 21968 31764 21974 31816
rect 22002 31764 22008 31816
rect 22060 31764 22066 31816
rect 22094 31764 22100 31816
rect 22152 31804 22158 31816
rect 22296 31813 22324 31844
rect 22189 31807 22247 31813
rect 22189 31804 22201 31807
rect 22152 31776 22201 31804
rect 22152 31764 22158 31776
rect 22189 31773 22201 31776
rect 22235 31773 22247 31807
rect 22189 31767 22247 31773
rect 22281 31807 22339 31813
rect 22281 31773 22293 31807
rect 22327 31773 22339 31807
rect 22281 31767 22339 31773
rect 22370 31764 22376 31816
rect 22428 31813 22434 31816
rect 22428 31804 22436 31813
rect 22649 31807 22707 31813
rect 22428 31776 22473 31804
rect 22428 31767 22436 31776
rect 22649 31773 22661 31807
rect 22695 31804 22707 31807
rect 22797 31807 22855 31813
rect 22695 31776 22729 31804
rect 22695 31773 22707 31776
rect 22649 31767 22707 31773
rect 22797 31773 22809 31807
rect 22843 31804 22855 31807
rect 22996 31804 23024 31844
rect 22843 31776 23024 31804
rect 22843 31773 22855 31776
rect 22797 31767 22855 31773
rect 22428 31764 22434 31767
rect 17218 31696 17224 31748
rect 17276 31736 17282 31748
rect 20530 31736 20536 31748
rect 17276 31708 20536 31736
rect 17276 31696 17282 31708
rect 20530 31696 20536 31708
rect 20588 31696 20594 31748
rect 22664 31680 22692 31767
rect 23106 31764 23112 31816
rect 23164 31813 23170 31816
rect 23164 31804 23172 31813
rect 23164 31776 23209 31804
rect 23164 31767 23172 31776
rect 23164 31764 23170 31767
rect 23290 31764 23296 31816
rect 23348 31804 23354 31816
rect 23492 31813 23520 31844
rect 23676 31844 24124 31872
rect 23676 31816 23704 31844
rect 24118 31832 24124 31844
rect 24176 31832 24182 31884
rect 23385 31807 23443 31813
rect 23385 31804 23397 31807
rect 23348 31776 23397 31804
rect 23348 31764 23354 31776
rect 23385 31773 23397 31776
rect 23431 31773 23443 31807
rect 23385 31767 23443 31773
rect 23478 31807 23536 31813
rect 23478 31773 23490 31807
rect 23524 31804 23536 31807
rect 23566 31804 23572 31816
rect 23524 31776 23572 31804
rect 23524 31773 23536 31776
rect 23478 31767 23536 31773
rect 23566 31764 23572 31776
rect 23624 31764 23630 31816
rect 23658 31764 23664 31816
rect 23716 31764 23722 31816
rect 23934 31813 23940 31816
rect 23891 31807 23940 31813
rect 23891 31773 23903 31807
rect 23937 31773 23940 31807
rect 23891 31767 23940 31773
rect 23934 31764 23940 31767
rect 23992 31804 23998 31816
rect 24210 31804 24216 31816
rect 23992 31776 24216 31804
rect 23992 31764 23998 31776
rect 24210 31764 24216 31776
rect 24268 31764 24274 31816
rect 24302 31764 24308 31816
rect 24360 31804 24366 31816
rect 24397 31807 24455 31813
rect 24397 31804 24409 31807
rect 24360 31776 24409 31804
rect 24360 31764 24366 31776
rect 24397 31773 24409 31776
rect 24443 31773 24455 31807
rect 24504 31804 24532 31912
rect 24949 31909 24961 31943
rect 24995 31909 25007 31943
rect 25056 31940 25084 31980
rect 25130 31968 25136 32020
rect 25188 32008 25194 32020
rect 32122 32008 32128 32020
rect 25188 31980 32128 32008
rect 25188 31968 25194 31980
rect 25225 31943 25283 31949
rect 25225 31940 25237 31943
rect 25056 31912 25237 31940
rect 24949 31903 25007 31909
rect 25225 31909 25237 31912
rect 25271 31909 25283 31943
rect 25225 31903 25283 31909
rect 24578 31832 24584 31884
rect 24636 31872 24642 31884
rect 24964 31872 24992 31903
rect 25498 31900 25504 31952
rect 25556 31940 25562 31952
rect 26789 31943 26847 31949
rect 26789 31940 26801 31943
rect 25556 31912 26801 31940
rect 25556 31900 25562 31912
rect 26789 31909 26801 31912
rect 26835 31909 26847 31943
rect 26789 31903 26847 31909
rect 26896 31872 26924 31980
rect 26970 31900 26976 31952
rect 27028 31900 27034 31952
rect 28718 31900 28724 31952
rect 28776 31940 28782 31952
rect 30193 31943 30251 31949
rect 28776 31912 29960 31940
rect 28776 31900 28782 31912
rect 24636 31844 24808 31872
rect 24964 31844 25452 31872
rect 24636 31832 24642 31844
rect 24780 31813 24808 31844
rect 24765 31807 24823 31813
rect 24504 31776 24716 31804
rect 24397 31767 24455 31773
rect 22922 31696 22928 31748
rect 22980 31696 22986 31748
rect 23017 31739 23075 31745
rect 23017 31705 23029 31739
rect 23063 31736 23075 31739
rect 23063 31708 23428 31736
rect 23063 31705 23075 31708
rect 23017 31699 23075 31705
rect 23400 31680 23428 31708
rect 23750 31696 23756 31748
rect 23808 31696 23814 31748
rect 24688 31745 24716 31776
rect 24765 31773 24777 31807
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 25038 31764 25044 31816
rect 25096 31764 25102 31816
rect 25130 31764 25136 31816
rect 25188 31764 25194 31816
rect 25314 31764 25320 31816
rect 25372 31764 25378 31816
rect 25424 31813 25452 31844
rect 26252 31844 26924 31872
rect 26988 31872 27016 31900
rect 29086 31872 29092 31884
rect 26988 31844 29092 31872
rect 25409 31807 25467 31813
rect 25409 31773 25421 31807
rect 25455 31773 25467 31807
rect 25409 31767 25467 31773
rect 26050 31764 26056 31816
rect 26108 31800 26114 31816
rect 26252 31813 26280 31844
rect 26145 31807 26203 31813
rect 26145 31800 26157 31807
rect 26108 31773 26157 31800
rect 26191 31773 26203 31807
rect 26108 31772 26203 31773
rect 26108 31764 26114 31772
rect 26145 31767 26203 31772
rect 26237 31807 26295 31813
rect 26237 31773 26249 31807
rect 26283 31773 26295 31807
rect 26237 31767 26295 31773
rect 26513 31807 26571 31813
rect 26513 31773 26525 31807
rect 26559 31804 26571 31807
rect 26694 31804 26700 31816
rect 26559 31776 26700 31804
rect 26559 31773 26571 31776
rect 26513 31767 26571 31773
rect 26694 31764 26700 31776
rect 26752 31764 26758 31816
rect 26988 31813 27016 31844
rect 29086 31832 29092 31844
rect 29144 31832 29150 31884
rect 26973 31807 27031 31813
rect 26973 31773 26985 31807
rect 27019 31773 27031 31807
rect 27890 31804 27896 31816
rect 26973 31767 27031 31773
rect 27356 31776 27896 31804
rect 24581 31739 24639 31745
rect 24581 31705 24593 31739
rect 24627 31705 24639 31739
rect 24581 31699 24639 31705
rect 24673 31739 24731 31745
rect 24673 31705 24685 31739
rect 24719 31736 24731 31739
rect 25056 31736 25084 31764
rect 27356 31748 27384 31776
rect 27890 31764 27896 31776
rect 27948 31804 27954 31816
rect 27985 31807 28043 31813
rect 27985 31804 27997 31807
rect 27948 31776 27997 31804
rect 27948 31764 27954 31776
rect 27985 31773 27997 31776
rect 28031 31773 28043 31807
rect 27985 31767 28043 31773
rect 28258 31764 28264 31816
rect 28316 31764 28322 31816
rect 29270 31764 29276 31816
rect 29328 31804 29334 31816
rect 29546 31804 29552 31816
rect 29328 31776 29552 31804
rect 29328 31764 29334 31776
rect 29546 31764 29552 31776
rect 29604 31764 29610 31816
rect 29642 31807 29700 31813
rect 29642 31773 29654 31807
rect 29688 31804 29700 31807
rect 29688 31776 29721 31804
rect 29688 31773 29700 31776
rect 29642 31767 29700 31773
rect 26329 31739 26387 31745
rect 26329 31736 26341 31739
rect 24719 31708 25084 31736
rect 25148 31708 26341 31736
rect 24719 31705 24731 31708
rect 24673 31699 24731 31705
rect 18138 31668 18144 31680
rect 16684 31640 18144 31668
rect 13449 31631 13507 31637
rect 18138 31628 18144 31640
rect 18196 31628 18202 31680
rect 18690 31628 18696 31680
rect 18748 31628 18754 31680
rect 19981 31671 20039 31677
rect 19981 31637 19993 31671
rect 20027 31668 20039 31671
rect 20162 31668 20168 31680
rect 20027 31640 20168 31668
rect 20027 31637 20039 31640
rect 19981 31631 20039 31637
rect 20162 31628 20168 31640
rect 20220 31628 20226 31680
rect 22554 31628 22560 31680
rect 22612 31628 22618 31680
rect 22646 31628 22652 31680
rect 22704 31628 22710 31680
rect 22738 31628 22744 31680
rect 22796 31668 22802 31680
rect 23293 31671 23351 31677
rect 23293 31668 23305 31671
rect 22796 31640 23305 31668
rect 22796 31628 22802 31640
rect 23293 31637 23305 31640
rect 23339 31637 23351 31671
rect 23293 31631 23351 31637
rect 23382 31628 23388 31680
rect 23440 31628 23446 31680
rect 24596 31668 24624 31699
rect 24762 31668 24768 31680
rect 24596 31640 24768 31668
rect 24762 31628 24768 31640
rect 24820 31628 24826 31680
rect 24946 31628 24952 31680
rect 25004 31668 25010 31680
rect 25148 31668 25176 31708
rect 25792 31680 25820 31708
rect 26329 31705 26341 31708
rect 26375 31705 26387 31739
rect 26329 31699 26387 31705
rect 27338 31696 27344 31748
rect 27396 31696 27402 31748
rect 25004 31640 25176 31668
rect 25004 31628 25010 31640
rect 25590 31628 25596 31680
rect 25648 31628 25654 31680
rect 25774 31628 25780 31680
rect 25832 31628 25838 31680
rect 25961 31671 26019 31677
rect 25961 31637 25973 31671
rect 26007 31668 26019 31671
rect 26142 31668 26148 31680
rect 26007 31640 26148 31668
rect 26007 31637 26019 31640
rect 25961 31631 26019 31637
rect 26142 31628 26148 31640
rect 26200 31628 26206 31680
rect 27706 31628 27712 31680
rect 27764 31668 27770 31680
rect 27893 31671 27951 31677
rect 27893 31668 27905 31671
rect 27764 31640 27905 31668
rect 27764 31628 27770 31640
rect 27893 31637 27905 31640
rect 27939 31637 27951 31671
rect 27893 31631 27951 31637
rect 27982 31628 27988 31680
rect 28040 31668 28046 31680
rect 28077 31671 28135 31677
rect 28077 31668 28089 31671
rect 28040 31640 28089 31668
rect 28040 31628 28046 31640
rect 28077 31637 28089 31640
rect 28123 31637 28135 31671
rect 28077 31631 28135 31637
rect 29546 31628 29552 31680
rect 29604 31668 29610 31680
rect 29656 31668 29684 31767
rect 29822 31764 29828 31816
rect 29880 31764 29886 31816
rect 29932 31813 29960 31912
rect 30193 31909 30205 31943
rect 30239 31940 30251 31943
rect 30239 31912 31800 31940
rect 30239 31909 30251 31912
rect 30193 31903 30251 31909
rect 30282 31832 30288 31884
rect 30340 31872 30346 31884
rect 30340 31844 30512 31872
rect 30340 31832 30346 31844
rect 29917 31807 29975 31813
rect 29917 31773 29929 31807
rect 29963 31773 29975 31807
rect 29917 31767 29975 31773
rect 30006 31764 30012 31816
rect 30064 31813 30070 31816
rect 30484 31813 30512 31844
rect 30064 31804 30072 31813
rect 30469 31807 30527 31813
rect 30064 31776 30157 31804
rect 30064 31767 30072 31776
rect 30469 31773 30481 31807
rect 30515 31773 30527 31807
rect 30469 31767 30527 31773
rect 30064 31764 30070 31767
rect 31478 31764 31484 31816
rect 31536 31764 31542 31816
rect 31772 31813 31800 31912
rect 31757 31807 31815 31813
rect 31757 31773 31769 31807
rect 31803 31773 31815 31807
rect 31757 31767 31815 31773
rect 30024 31736 30052 31764
rect 31573 31739 31631 31745
rect 30024 31708 30788 31736
rect 30760 31680 30788 31708
rect 31573 31705 31585 31739
rect 31619 31736 31631 31739
rect 31864 31736 31892 31980
rect 32122 31968 32128 31980
rect 32180 31968 32186 32020
rect 34606 31764 34612 31816
rect 34664 31804 34670 31816
rect 34885 31807 34943 31813
rect 34885 31804 34897 31807
rect 34664 31776 34897 31804
rect 34664 31764 34670 31776
rect 34885 31773 34897 31776
rect 34931 31804 34943 31807
rect 34977 31807 35035 31813
rect 34977 31804 34989 31807
rect 34931 31776 34989 31804
rect 34931 31773 34943 31776
rect 34885 31767 34943 31773
rect 34977 31773 34989 31776
rect 35023 31773 35035 31807
rect 34977 31767 35035 31773
rect 35434 31764 35440 31816
rect 35492 31764 35498 31816
rect 31619 31708 31892 31736
rect 31619 31705 31631 31708
rect 31573 31699 31631 31705
rect 34514 31696 34520 31748
rect 34572 31736 34578 31748
rect 35069 31739 35127 31745
rect 35069 31736 35081 31739
rect 34572 31708 35081 31736
rect 34572 31696 34578 31708
rect 35069 31705 35081 31708
rect 35115 31705 35127 31739
rect 35069 31699 35127 31705
rect 29604 31640 29684 31668
rect 29604 31628 29610 31640
rect 30374 31628 30380 31680
rect 30432 31628 30438 31680
rect 30742 31628 30748 31680
rect 30800 31628 30806 31680
rect 31941 31671 31999 31677
rect 31941 31637 31953 31671
rect 31987 31668 31999 31671
rect 32030 31668 32036 31680
rect 31987 31640 32036 31668
rect 31987 31637 31999 31640
rect 31941 31631 31999 31637
rect 32030 31628 32036 31640
rect 32088 31628 32094 31680
rect 34790 31628 34796 31680
rect 34848 31628 34854 31680
rect 35250 31628 35256 31680
rect 35308 31628 35314 31680
rect 1104 31578 38272 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38272 31578
rect 1104 31504 38272 31526
rect 8294 31464 8300 31476
rect 8128 31436 8300 31464
rect 8128 31405 8156 31436
rect 8294 31424 8300 31436
rect 8352 31424 8358 31476
rect 8938 31424 8944 31476
rect 8996 31464 9002 31476
rect 9490 31464 9496 31476
rect 8996 31436 9496 31464
rect 8996 31424 9002 31436
rect 9490 31424 9496 31436
rect 9548 31424 9554 31476
rect 9766 31424 9772 31476
rect 9824 31464 9830 31476
rect 9861 31467 9919 31473
rect 9861 31464 9873 31467
rect 9824 31436 9873 31464
rect 9824 31424 9830 31436
rect 9861 31433 9873 31436
rect 9907 31433 9919 31467
rect 9861 31427 9919 31433
rect 10137 31467 10195 31473
rect 10137 31433 10149 31467
rect 10183 31433 10195 31467
rect 10137 31427 10195 31433
rect 8113 31399 8171 31405
rect 8113 31365 8125 31399
rect 8159 31365 8171 31399
rect 8113 31359 8171 31365
rect 8386 31356 8392 31408
rect 8444 31396 8450 31408
rect 8444 31368 8602 31396
rect 8444 31356 8450 31368
rect 10045 31331 10103 31337
rect 10045 31297 10057 31331
rect 10091 31328 10103 31331
rect 10152 31328 10180 31427
rect 10502 31424 10508 31476
rect 10560 31464 10566 31476
rect 10962 31464 10968 31476
rect 10560 31436 10968 31464
rect 10560 31424 10566 31436
rect 10962 31424 10968 31436
rect 11020 31424 11026 31476
rect 13446 31424 13452 31476
rect 13504 31424 13510 31476
rect 16666 31464 16672 31476
rect 14660 31436 16672 31464
rect 11701 31399 11759 31405
rect 11701 31365 11713 31399
rect 11747 31396 11759 31399
rect 11974 31396 11980 31408
rect 11747 31368 11980 31396
rect 11747 31365 11759 31368
rect 11701 31359 11759 31365
rect 11974 31356 11980 31368
rect 12032 31396 12038 31408
rect 12526 31396 12532 31408
rect 12032 31368 12532 31396
rect 12032 31356 12038 31368
rect 12526 31356 12532 31368
rect 12584 31356 12590 31408
rect 14660 31396 14688 31436
rect 16666 31424 16672 31436
rect 16724 31424 16730 31476
rect 17313 31467 17371 31473
rect 17313 31433 17325 31467
rect 17359 31464 17371 31467
rect 18598 31464 18604 31476
rect 17359 31436 18604 31464
rect 17359 31433 17371 31436
rect 17313 31427 17371 31433
rect 18598 31424 18604 31436
rect 18656 31424 18662 31476
rect 18690 31424 18696 31476
rect 18748 31424 18754 31476
rect 21174 31424 21180 31476
rect 21232 31464 21238 31476
rect 21358 31464 21364 31476
rect 21232 31436 21364 31464
rect 21232 31424 21238 31436
rect 21358 31424 21364 31436
rect 21416 31424 21422 31476
rect 21450 31424 21456 31476
rect 21508 31464 21514 31476
rect 22097 31467 22155 31473
rect 22097 31464 22109 31467
rect 21508 31436 22109 31464
rect 21508 31424 21514 31436
rect 22097 31433 22109 31436
rect 22143 31433 22155 31467
rect 22097 31427 22155 31433
rect 22186 31424 22192 31476
rect 22244 31424 22250 31476
rect 22373 31467 22431 31473
rect 22373 31433 22385 31467
rect 22419 31464 22431 31467
rect 23290 31464 23296 31476
rect 22419 31436 23296 31464
rect 22419 31433 22431 31436
rect 22373 31427 22431 31433
rect 23290 31424 23296 31436
rect 23348 31424 23354 31476
rect 27614 31424 27620 31476
rect 27672 31424 27678 31476
rect 30374 31424 30380 31476
rect 30432 31424 30438 31476
rect 34790 31424 34796 31476
rect 34848 31424 34854 31476
rect 12912 31368 14688 31396
rect 14737 31399 14795 31405
rect 10091 31300 10180 31328
rect 10505 31331 10563 31337
rect 10091 31297 10103 31300
rect 10045 31291 10103 31297
rect 10505 31297 10517 31331
rect 10551 31328 10563 31331
rect 11517 31331 11575 31337
rect 11517 31328 11529 31331
rect 10551 31300 11529 31328
rect 10551 31297 10563 31300
rect 10505 31291 10563 31297
rect 11517 31297 11529 31300
rect 11563 31328 11575 31331
rect 11606 31328 11612 31340
rect 11563 31300 11612 31328
rect 11563 31297 11575 31300
rect 11517 31291 11575 31297
rect 11606 31288 11612 31300
rect 11664 31288 11670 31340
rect 11793 31331 11851 31337
rect 11793 31297 11805 31331
rect 11839 31297 11851 31331
rect 11793 31291 11851 31297
rect 7834 31220 7840 31272
rect 7892 31220 7898 31272
rect 10226 31220 10232 31272
rect 10284 31260 10290 31272
rect 10597 31263 10655 31269
rect 10597 31260 10609 31263
rect 10284 31232 10609 31260
rect 10284 31220 10290 31232
rect 10597 31229 10609 31232
rect 10643 31229 10655 31263
rect 10597 31223 10655 31229
rect 10781 31263 10839 31269
rect 10781 31229 10793 31263
rect 10827 31260 10839 31263
rect 10962 31260 10968 31272
rect 10827 31232 10968 31260
rect 10827 31229 10839 31232
rect 10781 31223 10839 31229
rect 10962 31220 10968 31232
rect 11020 31220 11026 31272
rect 11808 31260 11836 31291
rect 11882 31288 11888 31340
rect 11940 31328 11946 31340
rect 12342 31328 12348 31340
rect 11940 31300 12348 31328
rect 11940 31288 11946 31300
rect 12342 31288 12348 31300
rect 12400 31288 12406 31340
rect 12912 31272 12940 31368
rect 14737 31365 14749 31399
rect 14783 31396 14795 31399
rect 15838 31396 15844 31408
rect 14783 31368 15844 31396
rect 14783 31365 14795 31368
rect 14737 31359 14795 31365
rect 15838 31356 15844 31368
rect 15896 31356 15902 31408
rect 16114 31356 16120 31408
rect 16172 31356 16178 31408
rect 16390 31356 16396 31408
rect 16448 31356 16454 31408
rect 16960 31368 17540 31396
rect 15470 31288 15476 31340
rect 15528 31288 15534 31340
rect 15657 31331 15715 31337
rect 15657 31297 15669 31331
rect 15703 31328 15715 31331
rect 15746 31328 15752 31340
rect 15703 31300 15752 31328
rect 15703 31297 15715 31300
rect 15657 31291 15715 31297
rect 15746 31288 15752 31300
rect 15804 31288 15810 31340
rect 15933 31331 15991 31337
rect 15933 31297 15945 31331
rect 15979 31328 15991 31331
rect 16022 31328 16028 31340
rect 15979 31300 16028 31328
rect 15979 31297 15991 31300
rect 15933 31291 15991 31297
rect 16022 31288 16028 31300
rect 16080 31288 16086 31340
rect 16206 31288 16212 31340
rect 16264 31288 16270 31340
rect 16301 31331 16359 31337
rect 16301 31297 16313 31331
rect 16347 31328 16359 31331
rect 16408 31328 16436 31356
rect 16960 31337 16988 31368
rect 16658 31332 16716 31337
rect 16347 31300 16436 31328
rect 16500 31331 16716 31332
rect 16500 31304 16670 31331
rect 16347 31297 16359 31300
rect 16301 31291 16359 31297
rect 12894 31260 12900 31272
rect 11808 31232 12900 31260
rect 9582 31152 9588 31204
rect 9640 31192 9646 31204
rect 11808 31192 11836 31232
rect 12894 31220 12900 31232
rect 12952 31220 12958 31272
rect 15381 31263 15439 31269
rect 15381 31260 15393 31263
rect 14660 31232 15393 31260
rect 9640 31164 11836 31192
rect 9640 31152 9646 31164
rect 14660 31136 14688 31232
rect 15381 31229 15393 31232
rect 15427 31229 15439 31263
rect 15381 31223 15439 31229
rect 15841 31263 15899 31269
rect 15841 31229 15853 31263
rect 15887 31260 15899 31263
rect 16500 31260 16528 31304
rect 16658 31297 16670 31304
rect 16704 31297 16716 31331
rect 16658 31291 16716 31297
rect 16817 31331 16875 31337
rect 16817 31297 16829 31331
rect 16863 31328 16875 31331
rect 16945 31331 17003 31337
rect 16863 31297 16896 31328
rect 16817 31291 16896 31297
rect 16945 31297 16957 31331
rect 16991 31297 17003 31331
rect 16945 31291 17003 31297
rect 17037 31331 17095 31337
rect 17037 31297 17049 31331
rect 17083 31297 17095 31331
rect 17037 31291 17095 31297
rect 17153 31331 17211 31337
rect 17153 31297 17165 31331
rect 17199 31328 17211 31331
rect 17310 31328 17316 31340
rect 17199 31300 17316 31328
rect 17199 31297 17211 31300
rect 17153 31291 17211 31297
rect 15887 31232 16528 31260
rect 15887 31229 15899 31232
rect 15841 31223 15899 31229
rect 16206 31152 16212 31204
rect 16264 31192 16270 31204
rect 16264 31164 16620 31192
rect 16264 31152 16270 31164
rect 12069 31127 12127 31133
rect 12069 31093 12081 31127
rect 12115 31124 12127 31127
rect 13538 31124 13544 31136
rect 12115 31096 13544 31124
rect 12115 31093 12127 31096
rect 12069 31087 12127 31093
rect 13538 31084 13544 31096
rect 13596 31084 13602 31136
rect 14642 31084 14648 31136
rect 14700 31084 14706 31136
rect 16482 31084 16488 31136
rect 16540 31084 16546 31136
rect 16592 31124 16620 31164
rect 16666 31152 16672 31204
rect 16724 31192 16730 31204
rect 16868 31192 16896 31291
rect 16724 31164 16896 31192
rect 16724 31152 16730 31164
rect 17052 31124 17080 31291
rect 17310 31288 17316 31300
rect 17368 31288 17374 31340
rect 17405 31331 17463 31337
rect 17405 31297 17417 31331
rect 17451 31297 17463 31331
rect 17405 31291 17463 31297
rect 17218 31152 17224 31204
rect 17276 31192 17282 31204
rect 17420 31192 17448 31291
rect 17512 31260 17540 31368
rect 17862 31356 17868 31408
rect 17920 31396 17926 31408
rect 19978 31396 19984 31408
rect 17920 31368 19984 31396
rect 17920 31356 17926 31368
rect 19978 31356 19984 31368
rect 20036 31396 20042 31408
rect 23385 31399 23443 31405
rect 23385 31396 23397 31399
rect 20036 31368 23397 31396
rect 20036 31356 20042 31368
rect 23385 31365 23397 31368
rect 23431 31365 23443 31399
rect 23385 31359 23443 31365
rect 25133 31399 25191 31405
rect 25133 31365 25145 31399
rect 25179 31396 25191 31399
rect 25498 31396 25504 31408
rect 25179 31368 25504 31396
rect 25179 31365 25191 31368
rect 25133 31359 25191 31365
rect 25498 31356 25504 31368
rect 25556 31396 25562 31408
rect 27632 31396 27660 31424
rect 25556 31368 27660 31396
rect 25556 31356 25562 31368
rect 27982 31356 27988 31408
rect 28040 31356 28046 31408
rect 30392 31396 30420 31424
rect 34808 31396 34836 31424
rect 29932 31368 30420 31396
rect 34440 31368 34836 31396
rect 17586 31288 17592 31340
rect 17644 31288 17650 31340
rect 17678 31288 17684 31340
rect 17736 31288 17742 31340
rect 17770 31288 17776 31340
rect 17828 31288 17834 31340
rect 18046 31288 18052 31340
rect 18104 31288 18110 31340
rect 18509 31331 18567 31337
rect 18509 31297 18521 31331
rect 18555 31328 18567 31331
rect 18690 31328 18696 31340
rect 18555 31300 18696 31328
rect 18555 31297 18567 31300
rect 18509 31291 18567 31297
rect 18690 31288 18696 31300
rect 18748 31288 18754 31340
rect 18782 31288 18788 31340
rect 18840 31288 18846 31340
rect 19150 31288 19156 31340
rect 19208 31328 19214 31340
rect 19245 31331 19303 31337
rect 19245 31328 19257 31331
rect 19208 31300 19257 31328
rect 19208 31288 19214 31300
rect 19245 31297 19257 31300
rect 19291 31297 19303 31331
rect 19245 31291 19303 31297
rect 19521 31331 19579 31337
rect 19521 31297 19533 31331
rect 19567 31297 19579 31331
rect 19521 31291 19579 31297
rect 18064 31260 18092 31288
rect 17512 31232 19334 31260
rect 17276 31164 17448 31192
rect 17276 31152 17282 31164
rect 19306 31136 19334 31232
rect 19536 31204 19564 31291
rect 19702 31288 19708 31340
rect 19760 31288 19766 31340
rect 20530 31288 20536 31340
rect 20588 31288 20594 31340
rect 20622 31288 20628 31340
rect 20680 31288 20686 31340
rect 20714 31288 20720 31340
rect 20772 31328 20778 31340
rect 20809 31331 20867 31337
rect 20809 31328 20821 31331
rect 20772 31300 20821 31328
rect 20772 31288 20778 31300
rect 20809 31297 20821 31300
rect 20855 31297 20867 31331
rect 20809 31291 20867 31297
rect 20901 31331 20959 31337
rect 20901 31297 20913 31331
rect 20947 31328 20959 31331
rect 20947 31300 21036 31328
rect 20947 31297 20959 31300
rect 20901 31291 20959 31297
rect 21008 31269 21036 31300
rect 21082 31288 21088 31340
rect 21140 31328 21146 31340
rect 21361 31331 21419 31337
rect 21361 31328 21373 31331
rect 21140 31300 21373 31328
rect 21140 31288 21146 31300
rect 21361 31297 21373 31300
rect 21407 31297 21419 31331
rect 21361 31291 21419 31297
rect 21453 31331 21511 31337
rect 21453 31297 21465 31331
rect 21499 31297 21511 31331
rect 21453 31291 21511 31297
rect 20993 31263 21051 31269
rect 20993 31229 21005 31263
rect 21039 31229 21051 31263
rect 20993 31223 21051 31229
rect 21174 31220 21180 31272
rect 21232 31220 21238 31272
rect 21269 31263 21327 31269
rect 21269 31229 21281 31263
rect 21315 31229 21327 31263
rect 21468 31260 21496 31291
rect 21634 31288 21640 31340
rect 21692 31328 21698 31340
rect 21818 31328 21824 31340
rect 21692 31300 21824 31328
rect 21692 31288 21698 31300
rect 21818 31288 21824 31300
rect 21876 31288 21882 31340
rect 22005 31331 22063 31337
rect 22005 31297 22017 31331
rect 22051 31297 22063 31331
rect 22005 31291 22063 31297
rect 21726 31260 21732 31272
rect 21468 31232 21732 31260
rect 21269 31223 21327 31229
rect 19518 31152 19524 31204
rect 19576 31152 19582 31204
rect 21284 31192 21312 31223
rect 21726 31220 21732 31232
rect 21784 31220 21790 31272
rect 21450 31192 21456 31204
rect 21284 31164 21456 31192
rect 21450 31152 21456 31164
rect 21508 31152 21514 31204
rect 21542 31152 21548 31204
rect 21600 31192 21606 31204
rect 22020 31192 22048 31291
rect 22554 31288 22560 31340
rect 22612 31288 22618 31340
rect 22830 31288 22836 31340
rect 22888 31288 22894 31340
rect 23014 31288 23020 31340
rect 23072 31288 23078 31340
rect 23290 31288 23296 31340
rect 23348 31288 23354 31340
rect 25406 31288 25412 31340
rect 25464 31288 25470 31340
rect 25590 31288 25596 31340
rect 25648 31288 25654 31340
rect 26329 31331 26387 31337
rect 26329 31297 26341 31331
rect 26375 31326 26387 31331
rect 26375 31297 26389 31326
rect 26329 31291 26389 31297
rect 22572 31260 22600 31288
rect 22925 31263 22983 31269
rect 22925 31260 22937 31263
rect 22572 31232 22937 31260
rect 22925 31229 22937 31232
rect 22971 31229 22983 31263
rect 22925 31223 22983 31229
rect 23109 31263 23167 31269
rect 23109 31229 23121 31263
rect 23155 31260 23167 31263
rect 24578 31260 24584 31272
rect 23155 31232 24584 31260
rect 23155 31229 23167 31232
rect 23109 31223 23167 31229
rect 24578 31220 24584 31232
rect 24636 31220 24642 31272
rect 26053 31263 26111 31269
rect 26053 31229 26065 31263
rect 26099 31229 26111 31263
rect 26361 31260 26389 31291
rect 26418 31288 26424 31340
rect 26476 31328 26482 31340
rect 26973 31331 27031 31337
rect 26973 31328 26985 31331
rect 26476 31300 26985 31328
rect 26476 31288 26482 31300
rect 26973 31297 26985 31300
rect 27019 31297 27031 31331
rect 26973 31291 27031 31297
rect 27154 31288 27160 31340
rect 27212 31288 27218 31340
rect 27249 31331 27307 31337
rect 27249 31297 27261 31331
rect 27295 31297 27307 31331
rect 27249 31291 27307 31297
rect 27341 31331 27399 31337
rect 27341 31297 27353 31331
rect 27387 31328 27399 31331
rect 27387 31300 27476 31328
rect 29118 31300 29224 31328
rect 27387 31297 27399 31300
rect 27341 31291 27399 31297
rect 26510 31260 26516 31272
rect 26361 31232 26516 31260
rect 26053 31223 26111 31229
rect 26068 31192 26096 31223
rect 26510 31220 26516 31232
rect 26568 31220 26574 31272
rect 26786 31220 26792 31272
rect 26844 31260 26850 31272
rect 27264 31260 27292 31291
rect 26844 31232 27292 31260
rect 26844 31220 26850 31232
rect 21600 31164 22048 31192
rect 22572 31164 26096 31192
rect 21600 31152 21606 31164
rect 16592 31096 17080 31124
rect 17862 31084 17868 31136
rect 17920 31124 17926 31136
rect 17957 31127 18015 31133
rect 17957 31124 17969 31127
rect 17920 31096 17969 31124
rect 17920 31084 17926 31096
rect 17957 31093 17969 31096
rect 18003 31093 18015 31127
rect 17957 31087 18015 31093
rect 18322 31084 18328 31136
rect 18380 31084 18386 31136
rect 19306 31096 19340 31136
rect 19334 31084 19340 31096
rect 19392 31084 19398 31136
rect 20349 31127 20407 31133
rect 20349 31093 20361 31127
rect 20395 31124 20407 31127
rect 22572 31124 22600 31164
rect 26694 31152 26700 31204
rect 26752 31152 26758 31204
rect 27448 31136 27476 31300
rect 27706 31220 27712 31272
rect 27764 31220 27770 31272
rect 29196 31204 29224 31300
rect 29638 31288 29644 31340
rect 29696 31288 29702 31340
rect 29932 31337 29960 31368
rect 29917 31331 29975 31337
rect 29917 31297 29929 31331
rect 29963 31297 29975 31331
rect 29917 31291 29975 31297
rect 31220 31300 31326 31328
rect 30193 31263 30251 31269
rect 30193 31260 30205 31263
rect 29840 31232 30205 31260
rect 29178 31152 29184 31204
rect 29236 31192 29242 31204
rect 29840 31201 29868 31232
rect 30193 31229 30205 31232
rect 30239 31229 30251 31263
rect 30193 31223 30251 31229
rect 29825 31195 29883 31201
rect 29236 31164 29776 31192
rect 29236 31152 29242 31164
rect 20395 31096 22600 31124
rect 22649 31127 22707 31133
rect 20395 31093 20407 31096
rect 20349 31087 20407 31093
rect 22649 31093 22661 31127
rect 22695 31124 22707 31127
rect 23014 31124 23020 31136
rect 22695 31096 23020 31124
rect 22695 31093 22707 31096
rect 22649 31087 22707 31093
rect 23014 31084 23020 31096
rect 23072 31084 23078 31136
rect 25406 31084 25412 31136
rect 25464 31124 25470 31136
rect 26418 31124 26424 31136
rect 25464 31096 26424 31124
rect 25464 31084 25470 31096
rect 26418 31084 26424 31096
rect 26476 31084 26482 31136
rect 27430 31084 27436 31136
rect 27488 31084 27494 31136
rect 27617 31127 27675 31133
rect 27617 31093 27629 31127
rect 27663 31124 27675 31127
rect 27706 31124 27712 31136
rect 27663 31096 27712 31124
rect 27663 31093 27675 31096
rect 27617 31087 27675 31093
rect 27706 31084 27712 31096
rect 27764 31084 27770 31136
rect 28994 31084 29000 31136
rect 29052 31124 29058 31136
rect 29457 31127 29515 31133
rect 29457 31124 29469 31127
rect 29052 31096 29469 31124
rect 29052 31084 29058 31096
rect 29457 31093 29469 31096
rect 29503 31124 29515 31127
rect 29546 31124 29552 31136
rect 29503 31096 29552 31124
rect 29503 31093 29515 31096
rect 29457 31087 29515 31093
rect 29546 31084 29552 31096
rect 29604 31084 29610 31136
rect 29748 31124 29776 31164
rect 29825 31161 29837 31195
rect 29871 31161 29883 31195
rect 29825 31155 29883 31161
rect 31220 31124 31248 31300
rect 31662 31288 31668 31340
rect 31720 31328 31726 31340
rect 34440 31337 34468 31368
rect 32401 31331 32459 31337
rect 32401 31328 32413 31331
rect 31720 31300 32413 31328
rect 31720 31288 31726 31300
rect 32401 31297 32413 31300
rect 32447 31297 32459 31331
rect 34425 31331 34483 31337
rect 32401 31291 32459 31297
rect 32968 31300 33074 31328
rect 31938 31220 31944 31272
rect 31996 31220 32002 31272
rect 32968 31136 32996 31300
rect 34425 31297 34437 31331
rect 34471 31297 34483 31331
rect 34425 31291 34483 31297
rect 34514 31288 34520 31340
rect 34572 31288 34578 31340
rect 35926 31300 36032 31328
rect 34146 31220 34152 31272
rect 34204 31220 34210 31272
rect 34793 31263 34851 31269
rect 34793 31229 34805 31263
rect 34839 31260 34851 31263
rect 35250 31260 35256 31272
rect 34839 31232 35256 31260
rect 34839 31229 34851 31232
rect 34793 31223 34851 31229
rect 35250 31220 35256 31232
rect 35308 31220 35314 31272
rect 36004 31136 36032 31300
rect 36538 31220 36544 31272
rect 36596 31220 36602 31272
rect 29748 31096 31248 31124
rect 32950 31084 32956 31136
rect 33008 31084 33014 31136
rect 35986 31084 35992 31136
rect 36044 31084 36050 31136
rect 1104 31034 38272 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38272 31034
rect 1104 30960 38272 30982
rect 6362 30880 6368 30932
rect 6420 30920 6426 30932
rect 8386 30920 8392 30932
rect 6420 30892 8392 30920
rect 6420 30880 6426 30892
rect 3970 30676 3976 30728
rect 4028 30716 4034 30728
rect 4525 30719 4583 30725
rect 4525 30716 4537 30719
rect 4028 30688 4537 30716
rect 4028 30676 4034 30688
rect 4525 30685 4537 30688
rect 4571 30685 4583 30719
rect 4525 30679 4583 30685
rect 5626 30676 5632 30728
rect 5684 30676 5690 30728
rect 5721 30719 5779 30725
rect 5721 30685 5733 30719
rect 5767 30716 5779 30719
rect 5905 30719 5963 30725
rect 5905 30716 5917 30719
rect 5767 30688 5917 30716
rect 5767 30685 5779 30688
rect 5721 30679 5779 30685
rect 5905 30685 5917 30688
rect 5951 30685 5963 30719
rect 7300 30702 7328 30892
rect 8386 30880 8392 30892
rect 8444 30880 8450 30932
rect 8478 30880 8484 30932
rect 8536 30920 8542 30932
rect 8941 30923 8999 30929
rect 8941 30920 8953 30923
rect 8536 30892 8953 30920
rect 8536 30880 8542 30892
rect 8941 30889 8953 30892
rect 8987 30889 8999 30923
rect 9582 30920 9588 30932
rect 8941 30883 8999 30889
rect 9416 30892 9588 30920
rect 7484 30824 8432 30852
rect 7484 30796 7512 30824
rect 7466 30744 7472 30796
rect 7524 30744 7530 30796
rect 8404 30793 8432 30824
rect 9416 30793 9444 30892
rect 9582 30880 9588 30892
rect 9640 30880 9646 30932
rect 14458 30880 14464 30932
rect 14516 30880 14522 30932
rect 16206 30880 16212 30932
rect 16264 30880 16270 30932
rect 16485 30923 16543 30929
rect 16485 30889 16497 30923
rect 16531 30920 16543 30923
rect 17586 30920 17592 30932
rect 16531 30892 17592 30920
rect 16531 30889 16543 30892
rect 16485 30883 16543 30889
rect 17586 30880 17592 30892
rect 17644 30880 17650 30932
rect 20990 30920 20996 30932
rect 18064 30892 20996 30920
rect 11606 30812 11612 30864
rect 11664 30852 11670 30864
rect 13357 30855 13415 30861
rect 13357 30852 13369 30855
rect 11664 30824 13369 30852
rect 11664 30812 11670 30824
rect 13357 30821 13369 30824
rect 13403 30852 13415 30855
rect 16224 30852 16252 30880
rect 18064 30864 18092 30892
rect 20990 30880 20996 30892
rect 21048 30880 21054 30932
rect 21269 30923 21327 30929
rect 21269 30889 21281 30923
rect 21315 30920 21327 30923
rect 21910 30920 21916 30932
rect 21315 30892 21916 30920
rect 21315 30889 21327 30892
rect 21269 30883 21327 30889
rect 21910 30880 21916 30892
rect 21968 30880 21974 30932
rect 24394 30880 24400 30932
rect 24452 30920 24458 30932
rect 24489 30923 24547 30929
rect 24489 30920 24501 30923
rect 24452 30892 24501 30920
rect 24452 30880 24458 30892
rect 24489 30889 24501 30892
rect 24535 30889 24547 30923
rect 24489 30883 24547 30889
rect 24857 30923 24915 30929
rect 24857 30889 24869 30923
rect 24903 30920 24915 30923
rect 25130 30920 25136 30932
rect 24903 30892 25136 30920
rect 24903 30889 24915 30892
rect 24857 30883 24915 30889
rect 25130 30880 25136 30892
rect 25188 30880 25194 30932
rect 26605 30923 26663 30929
rect 25976 30892 26556 30920
rect 13403 30824 16252 30852
rect 13403 30821 13415 30824
rect 13357 30815 13415 30821
rect 16850 30812 16856 30864
rect 16908 30852 16914 30864
rect 17126 30852 17132 30864
rect 16908 30824 17132 30852
rect 16908 30812 16914 30824
rect 17126 30812 17132 30824
rect 17184 30812 17190 30864
rect 18046 30812 18052 30864
rect 18104 30812 18110 30864
rect 20346 30812 20352 30864
rect 20404 30812 20410 30864
rect 20714 30812 20720 30864
rect 20772 30812 20778 30864
rect 21008 30852 21036 30880
rect 21729 30855 21787 30861
rect 21729 30852 21741 30855
rect 21008 30824 21741 30852
rect 21729 30821 21741 30824
rect 21775 30852 21787 30855
rect 22554 30852 22560 30864
rect 21775 30824 22560 30852
rect 21775 30821 21787 30824
rect 21729 30815 21787 30821
rect 22554 30812 22560 30824
rect 22612 30852 22618 30864
rect 23290 30852 23296 30864
rect 22612 30824 23296 30852
rect 22612 30812 22618 30824
rect 23290 30812 23296 30824
rect 23348 30812 23354 30864
rect 7653 30787 7711 30793
rect 7653 30753 7665 30787
rect 7699 30784 7711 30787
rect 8389 30787 8447 30793
rect 7699 30756 8248 30784
rect 7699 30753 7711 30756
rect 7653 30747 7711 30753
rect 8220 30725 8248 30756
rect 8389 30753 8401 30787
rect 8435 30753 8447 30787
rect 8389 30747 8447 30753
rect 9401 30787 9459 30793
rect 9401 30753 9413 30787
rect 9447 30753 9459 30787
rect 9401 30747 9459 30753
rect 9490 30744 9496 30796
rect 9548 30744 9554 30796
rect 13909 30787 13967 30793
rect 13909 30753 13921 30787
rect 13955 30784 13967 30787
rect 14553 30787 14611 30793
rect 14553 30784 14565 30787
rect 13955 30756 14565 30784
rect 13955 30753 13967 30756
rect 13909 30747 13967 30753
rect 14553 30753 14565 30756
rect 14599 30753 14611 30787
rect 14553 30747 14611 30753
rect 16942 30744 16948 30796
rect 17000 30784 17006 30796
rect 24578 30784 24584 30796
rect 17000 30756 24584 30784
rect 17000 30744 17006 30756
rect 24578 30744 24584 30756
rect 24636 30784 24642 30796
rect 25976 30784 26004 30892
rect 26528 30852 26556 30892
rect 26605 30889 26617 30923
rect 26651 30920 26663 30923
rect 27154 30920 27160 30932
rect 26651 30892 27160 30920
rect 26651 30889 26663 30892
rect 26605 30883 26663 30889
rect 27154 30880 27160 30892
rect 27212 30880 27218 30932
rect 28077 30923 28135 30929
rect 28077 30889 28089 30923
rect 28123 30920 28135 30923
rect 28258 30920 28264 30932
rect 28123 30892 28264 30920
rect 28123 30889 28135 30892
rect 28077 30883 28135 30889
rect 28258 30880 28264 30892
rect 28316 30880 28322 30932
rect 29638 30880 29644 30932
rect 29696 30920 29702 30932
rect 30101 30923 30159 30929
rect 30101 30920 30113 30923
rect 29696 30892 30113 30920
rect 29696 30880 29702 30892
rect 30101 30889 30113 30892
rect 30147 30889 30159 30923
rect 30101 30883 30159 30889
rect 33318 30880 33324 30932
rect 33376 30920 33382 30932
rect 34057 30923 34115 30929
rect 33376 30892 34008 30920
rect 33376 30880 33382 30892
rect 33781 30855 33839 30861
rect 26528 30824 27476 30852
rect 26786 30784 26792 30796
rect 24636 30756 26004 30784
rect 26252 30756 26792 30784
rect 24636 30744 24642 30756
rect 8205 30719 8263 30725
rect 5905 30679 5963 30685
rect 8205 30685 8217 30719
rect 8251 30716 8263 30719
rect 11698 30716 11704 30728
rect 8251 30688 11704 30716
rect 8251 30685 8263 30688
rect 8205 30679 8263 30685
rect 11698 30676 11704 30688
rect 11756 30716 11762 30728
rect 14369 30719 14427 30725
rect 11756 30688 14320 30716
rect 11756 30676 11762 30688
rect 4246 30540 4252 30592
rect 4304 30580 4310 30592
rect 4433 30583 4491 30589
rect 4433 30580 4445 30583
rect 4304 30552 4445 30580
rect 4304 30540 4310 30552
rect 4433 30549 4445 30552
rect 4479 30549 4491 30583
rect 5644 30580 5672 30676
rect 6178 30608 6184 30660
rect 6236 30608 6242 30660
rect 9582 30648 9588 30660
rect 7484 30620 9588 30648
rect 7484 30580 7512 30620
rect 9582 30608 9588 30620
rect 9640 30608 9646 30660
rect 13262 30608 13268 30660
rect 13320 30608 13326 30660
rect 13354 30608 13360 30660
rect 13412 30648 13418 30660
rect 13412 30620 13676 30648
rect 13412 30608 13418 30620
rect 5644 30552 7512 30580
rect 4433 30543 4491 30549
rect 7834 30540 7840 30592
rect 7892 30540 7898 30592
rect 8018 30540 8024 30592
rect 8076 30580 8082 30592
rect 8297 30583 8355 30589
rect 8297 30580 8309 30583
rect 8076 30552 8309 30580
rect 8076 30540 8082 30552
rect 8297 30549 8309 30552
rect 8343 30580 8355 30583
rect 9309 30583 9367 30589
rect 9309 30580 9321 30583
rect 8343 30552 9321 30580
rect 8343 30549 8355 30552
rect 8297 30543 8355 30549
rect 9309 30549 9321 30552
rect 9355 30580 9367 30583
rect 10226 30580 10232 30592
rect 9355 30552 10232 30580
rect 9355 30549 9367 30552
rect 9309 30543 9367 30549
rect 10226 30540 10232 30552
rect 10284 30540 10290 30592
rect 13280 30580 13308 30608
rect 13648 30589 13676 30620
rect 13722 30608 13728 30660
rect 13780 30608 13786 30660
rect 14292 30648 14320 30688
rect 14369 30685 14381 30719
rect 14415 30716 14427 30719
rect 14458 30716 14464 30728
rect 14415 30688 14464 30716
rect 14415 30685 14427 30688
rect 14369 30679 14427 30685
rect 14458 30676 14464 30688
rect 14516 30676 14522 30728
rect 14642 30676 14648 30728
rect 14700 30676 14706 30728
rect 14734 30676 14740 30728
rect 14792 30716 14798 30728
rect 14829 30719 14887 30725
rect 14829 30716 14841 30719
rect 14792 30688 14841 30716
rect 14792 30676 14798 30688
rect 14829 30685 14841 30688
rect 14875 30685 14887 30719
rect 16301 30719 16359 30725
rect 16301 30716 16313 30719
rect 14829 30679 14887 30685
rect 14936 30688 16313 30716
rect 14660 30648 14688 30676
rect 14936 30648 14964 30688
rect 16301 30685 16313 30688
rect 16347 30685 16359 30719
rect 16301 30679 16359 30685
rect 16574 30676 16580 30728
rect 16632 30676 16638 30728
rect 16666 30676 16672 30728
rect 16724 30716 16730 30728
rect 16724 30688 16769 30716
rect 16724 30676 16730 30688
rect 16850 30676 16856 30728
rect 16908 30676 16914 30728
rect 17083 30719 17141 30725
rect 17083 30685 17095 30719
rect 17129 30716 17141 30719
rect 17402 30716 17408 30728
rect 17129 30688 17408 30716
rect 17129 30685 17141 30688
rect 17083 30679 17141 30685
rect 17402 30676 17408 30688
rect 17460 30716 17466 30728
rect 17586 30716 17592 30728
rect 17460 30688 17592 30716
rect 17460 30676 17466 30688
rect 17586 30676 17592 30688
rect 17644 30676 17650 30728
rect 19058 30676 19064 30728
rect 19116 30676 19122 30728
rect 19518 30676 19524 30728
rect 19576 30676 19582 30728
rect 20254 30676 20260 30728
rect 20312 30676 20318 30728
rect 20438 30676 20444 30728
rect 20496 30716 20502 30728
rect 21085 30719 21143 30725
rect 20496 30688 21036 30716
rect 20496 30676 20502 30688
rect 14016 30620 14228 30648
rect 14292 30620 14964 30648
rect 16117 30651 16175 30657
rect 13541 30583 13599 30589
rect 13541 30580 13553 30583
rect 13280 30552 13553 30580
rect 13541 30549 13553 30552
rect 13587 30549 13599 30583
rect 13541 30543 13599 30549
rect 13633 30583 13691 30589
rect 13633 30549 13645 30583
rect 13679 30580 13691 30583
rect 14016 30580 14044 30620
rect 13679 30552 14044 30580
rect 13679 30549 13691 30552
rect 13633 30543 13691 30549
rect 14090 30540 14096 30592
rect 14148 30540 14154 30592
rect 14200 30580 14228 30620
rect 16117 30617 16129 30651
rect 16163 30617 16175 30651
rect 16117 30611 16175 30617
rect 16945 30651 17003 30657
rect 16945 30617 16957 30651
rect 16991 30617 17003 30651
rect 16945 30611 17003 30617
rect 14366 30580 14372 30592
rect 14200 30552 14372 30580
rect 14366 30540 14372 30552
rect 14424 30540 14430 30592
rect 15930 30540 15936 30592
rect 15988 30580 15994 30592
rect 16132 30580 16160 30611
rect 16298 30580 16304 30592
rect 15988 30552 16304 30580
rect 15988 30540 15994 30552
rect 16298 30540 16304 30552
rect 16356 30540 16362 30592
rect 16666 30540 16672 30592
rect 16724 30580 16730 30592
rect 16960 30580 16988 30611
rect 18506 30608 18512 30660
rect 18564 30648 18570 30660
rect 20346 30648 20352 30660
rect 18564 30620 20352 30648
rect 18564 30608 18570 30620
rect 20346 30608 20352 30620
rect 20404 30608 20410 30660
rect 21008 30657 21036 30688
rect 21085 30685 21097 30719
rect 21131 30716 21143 30719
rect 21266 30716 21272 30728
rect 21131 30688 21272 30716
rect 21131 30685 21143 30688
rect 21085 30679 21143 30685
rect 21266 30676 21272 30688
rect 21324 30676 21330 30728
rect 21358 30676 21364 30728
rect 21416 30676 21422 30728
rect 24489 30719 24547 30725
rect 24489 30685 24501 30719
rect 24535 30685 24547 30719
rect 24489 30679 24547 30685
rect 20993 30651 21051 30657
rect 20993 30617 21005 30651
rect 21039 30617 21051 30651
rect 21284 30648 21312 30676
rect 21545 30651 21603 30657
rect 21545 30648 21557 30651
rect 21284 30620 21557 30648
rect 20993 30611 21051 30617
rect 21545 30617 21557 30620
rect 21591 30617 21603 30651
rect 24504 30648 24532 30679
rect 25406 30676 25412 30728
rect 25464 30716 25470 30728
rect 25958 30716 25964 30728
rect 25464 30688 25964 30716
rect 25464 30676 25470 30688
rect 25958 30676 25964 30688
rect 26016 30716 26022 30728
rect 26053 30719 26111 30725
rect 26053 30716 26065 30719
rect 26016 30688 26065 30716
rect 26016 30676 26022 30688
rect 26053 30685 26065 30688
rect 26099 30685 26111 30719
rect 26053 30679 26111 30685
rect 26142 30676 26148 30728
rect 26200 30676 26206 30728
rect 24578 30648 24584 30660
rect 24504 30620 24584 30648
rect 21545 30611 21603 30617
rect 24578 30608 24584 30620
rect 24636 30648 24642 30660
rect 26252 30648 26280 30756
rect 26786 30744 26792 30756
rect 26844 30744 26850 30796
rect 27448 30728 27476 30824
rect 33781 30821 33793 30855
rect 33827 30821 33839 30855
rect 33781 30815 33839 30821
rect 27614 30744 27620 30796
rect 27672 30784 27678 30796
rect 28626 30784 28632 30796
rect 27672 30756 28632 30784
rect 27672 30744 27678 30756
rect 28626 30744 28632 30756
rect 28684 30744 28690 30796
rect 30650 30744 30656 30796
rect 30708 30744 30714 30796
rect 31018 30744 31024 30796
rect 31076 30784 31082 30796
rect 31662 30784 31668 30796
rect 31076 30756 31668 30784
rect 31076 30744 31082 30756
rect 31662 30744 31668 30756
rect 31720 30784 31726 30796
rect 31720 30756 32628 30784
rect 31720 30744 31726 30756
rect 26329 30719 26387 30725
rect 26329 30685 26341 30719
rect 26375 30685 26387 30719
rect 26329 30679 26387 30685
rect 24636 30620 26280 30648
rect 26344 30648 26372 30679
rect 26418 30676 26424 30728
rect 26476 30716 26482 30728
rect 26602 30716 26608 30728
rect 26476 30688 26608 30716
rect 26476 30676 26482 30688
rect 26602 30676 26608 30688
rect 26660 30676 26666 30728
rect 27430 30676 27436 30728
rect 27488 30716 27494 30728
rect 30469 30719 30527 30725
rect 30469 30716 30481 30719
rect 27488 30688 30481 30716
rect 27488 30676 27494 30688
rect 30469 30685 30481 30688
rect 30515 30716 30527 30719
rect 31938 30716 31944 30728
rect 30515 30688 31944 30716
rect 30515 30685 30527 30688
rect 30469 30679 30527 30685
rect 31938 30676 31944 30688
rect 31996 30716 32002 30728
rect 32490 30716 32496 30728
rect 31996 30688 32496 30716
rect 31996 30676 32002 30688
rect 32490 30676 32496 30688
rect 32548 30676 32554 30728
rect 32600 30716 32628 30756
rect 32766 30744 32772 30796
rect 32824 30784 32830 30796
rect 33134 30784 33140 30796
rect 32824 30756 33140 30784
rect 32824 30744 32830 30756
rect 33134 30744 33140 30756
rect 33192 30744 33198 30796
rect 33413 30719 33471 30725
rect 33413 30716 33425 30719
rect 32600 30688 33425 30716
rect 33413 30685 33425 30688
rect 33459 30685 33471 30719
rect 33796 30716 33824 30815
rect 33980 30796 34008 30892
rect 34057 30889 34069 30923
rect 34103 30920 34115 30923
rect 34146 30920 34152 30932
rect 34103 30892 34152 30920
rect 34103 30889 34115 30892
rect 34057 30883 34115 30889
rect 34146 30880 34152 30892
rect 34204 30880 34210 30932
rect 35434 30880 35440 30932
rect 35492 30880 35498 30932
rect 33962 30744 33968 30796
rect 34020 30784 34026 30796
rect 34793 30787 34851 30793
rect 34793 30784 34805 30787
rect 34020 30756 34805 30784
rect 34020 30744 34026 30756
rect 34793 30753 34805 30756
rect 34839 30753 34851 30787
rect 34793 30747 34851 30753
rect 33873 30719 33931 30725
rect 33873 30716 33885 30719
rect 33796 30688 33885 30716
rect 33413 30679 33471 30685
rect 33873 30685 33885 30688
rect 33919 30685 33931 30719
rect 33873 30679 33931 30685
rect 28537 30651 28595 30657
rect 28537 30648 28549 30651
rect 26344 30620 28549 30648
rect 24636 30608 24642 30620
rect 16724 30552 16988 30580
rect 16724 30540 16730 30552
rect 17218 30540 17224 30592
rect 17276 30540 17282 30592
rect 17773 30583 17831 30589
rect 17773 30549 17785 30583
rect 17819 30580 17831 30583
rect 17954 30580 17960 30592
rect 17819 30552 17960 30580
rect 17819 30549 17831 30552
rect 17773 30543 17831 30549
rect 17954 30540 17960 30552
rect 18012 30540 18018 30592
rect 18138 30540 18144 30592
rect 18196 30580 18202 30592
rect 18782 30580 18788 30592
rect 18196 30552 18788 30580
rect 18196 30540 18202 30552
rect 18782 30540 18788 30552
rect 18840 30580 18846 30592
rect 19518 30580 19524 30592
rect 18840 30552 19524 30580
rect 18840 30540 18846 30552
rect 19518 30540 19524 30552
rect 19576 30540 19582 30592
rect 20070 30540 20076 30592
rect 20128 30580 20134 30592
rect 20898 30580 20904 30592
rect 20128 30552 20904 30580
rect 20128 30540 20134 30552
rect 20898 30540 20904 30552
rect 20956 30540 20962 30592
rect 23566 30540 23572 30592
rect 23624 30580 23630 30592
rect 26344 30580 26372 30620
rect 28537 30617 28549 30620
rect 28583 30648 28595 30651
rect 28994 30648 29000 30660
rect 28583 30620 29000 30648
rect 28583 30617 28595 30620
rect 28537 30611 28595 30617
rect 28994 30608 29000 30620
rect 29052 30608 29058 30660
rect 30926 30608 30932 30660
rect 30984 30608 30990 30660
rect 33686 30608 33692 30660
rect 33744 30648 33750 30660
rect 34977 30651 35035 30657
rect 34977 30648 34989 30651
rect 33744 30620 34989 30648
rect 33744 30608 33750 30620
rect 34977 30617 34989 30620
rect 35023 30648 35035 30651
rect 36538 30648 36544 30660
rect 35023 30620 36544 30648
rect 35023 30617 35035 30620
rect 34977 30611 35035 30617
rect 36538 30608 36544 30620
rect 36596 30608 36602 30660
rect 23624 30552 26372 30580
rect 23624 30540 23630 30552
rect 28442 30540 28448 30592
rect 28500 30580 28506 30592
rect 30561 30583 30619 30589
rect 30561 30580 30573 30583
rect 28500 30552 30573 30580
rect 28500 30540 28506 30552
rect 30561 30549 30573 30552
rect 30607 30580 30619 30583
rect 30834 30580 30840 30592
rect 30607 30552 30840 30580
rect 30607 30549 30619 30552
rect 30561 30543 30619 30549
rect 30834 30540 30840 30552
rect 30892 30540 30898 30592
rect 31294 30540 31300 30592
rect 31352 30580 31358 30592
rect 32217 30583 32275 30589
rect 32217 30580 32229 30583
rect 31352 30552 32229 30580
rect 31352 30540 31358 30552
rect 32217 30549 32229 30552
rect 32263 30549 32275 30583
rect 32217 30543 32275 30549
rect 33318 30540 33324 30592
rect 33376 30580 33382 30592
rect 35069 30583 35127 30589
rect 35069 30580 35081 30583
rect 33376 30552 35081 30580
rect 33376 30540 33382 30552
rect 35069 30549 35081 30552
rect 35115 30549 35127 30583
rect 35069 30543 35127 30549
rect 1104 30490 38272 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38272 30490
rect 1104 30416 38272 30438
rect 5997 30379 6055 30385
rect 5997 30345 6009 30379
rect 6043 30345 6055 30379
rect 5997 30339 6055 30345
rect 5258 30268 5264 30320
rect 5316 30268 5322 30320
rect 6012 30240 6040 30339
rect 6178 30336 6184 30388
rect 6236 30376 6242 30388
rect 6457 30379 6515 30385
rect 6457 30376 6469 30379
rect 6236 30348 6469 30376
rect 6236 30336 6242 30348
rect 6457 30345 6469 30348
rect 6503 30345 6515 30379
rect 7650 30376 7656 30388
rect 6457 30339 6515 30345
rect 7208 30348 7656 30376
rect 6641 30243 6699 30249
rect 6012 30212 6592 30240
rect 4246 30132 4252 30184
rect 4304 30132 4310 30184
rect 4525 30175 4583 30181
rect 4525 30141 4537 30175
rect 4571 30172 4583 30175
rect 6564 30172 6592 30212
rect 6641 30209 6653 30243
rect 6687 30240 6699 30243
rect 7208 30240 7236 30348
rect 7650 30336 7656 30348
rect 7708 30336 7714 30388
rect 7742 30336 7748 30388
rect 7800 30376 7806 30388
rect 8018 30376 8024 30388
rect 7800 30348 8024 30376
rect 7800 30336 7806 30348
rect 8018 30336 8024 30348
rect 8076 30336 8082 30388
rect 9582 30336 9588 30388
rect 9640 30376 9646 30388
rect 13446 30376 13452 30388
rect 9640 30348 13452 30376
rect 9640 30336 9646 30348
rect 13446 30336 13452 30348
rect 13504 30336 13510 30388
rect 15010 30336 15016 30388
rect 15068 30376 15074 30388
rect 18046 30376 18052 30388
rect 15068 30348 18052 30376
rect 15068 30336 15074 30348
rect 18046 30336 18052 30348
rect 18104 30336 18110 30388
rect 19794 30336 19800 30388
rect 19852 30376 19858 30388
rect 20257 30379 20315 30385
rect 19852 30348 20116 30376
rect 19852 30336 19858 30348
rect 7377 30311 7435 30317
rect 7377 30277 7389 30311
rect 7423 30308 7435 30311
rect 7423 30280 8064 30308
rect 7423 30277 7435 30280
rect 7377 30271 7435 30277
rect 6687 30212 7236 30240
rect 6687 30209 6699 30212
rect 6641 30203 6699 30209
rect 7282 30200 7288 30252
rect 7340 30240 7346 30252
rect 7653 30243 7711 30249
rect 7653 30240 7665 30243
rect 7340 30212 7665 30240
rect 7340 30200 7346 30212
rect 7653 30209 7665 30212
rect 7699 30209 7711 30243
rect 7653 30203 7711 30209
rect 7742 30200 7748 30252
rect 7800 30200 7806 30252
rect 7837 30243 7895 30249
rect 7837 30209 7849 30243
rect 7883 30240 7895 30243
rect 7926 30240 7932 30252
rect 7883 30212 7932 30240
rect 7883 30209 7895 30212
rect 7837 30203 7895 30209
rect 7926 30200 7932 30212
rect 7984 30200 7990 30252
rect 8036 30249 8064 30280
rect 9950 30268 9956 30320
rect 10008 30308 10014 30320
rect 12989 30311 13047 30317
rect 12989 30308 13001 30311
rect 10008 30280 13001 30308
rect 10008 30268 10014 30280
rect 12989 30277 13001 30280
rect 13035 30277 13047 30311
rect 12989 30271 13047 30277
rect 14737 30311 14795 30317
rect 14737 30277 14749 30311
rect 14783 30308 14795 30311
rect 19518 30308 19524 30320
rect 14783 30280 19524 30308
rect 14783 30277 14795 30280
rect 14737 30271 14795 30277
rect 19518 30268 19524 30280
rect 19576 30268 19582 30320
rect 19889 30311 19947 30317
rect 19889 30277 19901 30311
rect 19935 30308 19947 30311
rect 19978 30308 19984 30320
rect 19935 30280 19984 30308
rect 19935 30277 19947 30280
rect 19889 30271 19947 30277
rect 8021 30243 8079 30249
rect 8021 30209 8033 30243
rect 8067 30209 8079 30243
rect 8021 30203 8079 30209
rect 8570 30200 8576 30252
rect 8628 30200 8634 30252
rect 9490 30200 9496 30252
rect 9548 30240 9554 30252
rect 10042 30240 10048 30252
rect 9548 30212 10048 30240
rect 9548 30200 9554 30212
rect 10042 30200 10048 30212
rect 10100 30200 10106 30252
rect 11514 30200 11520 30252
rect 11572 30240 11578 30252
rect 11609 30243 11667 30249
rect 11609 30240 11621 30243
rect 11572 30212 11621 30240
rect 11572 30200 11578 30212
rect 11609 30209 11621 30212
rect 11655 30209 11667 30243
rect 11609 30203 11667 30209
rect 11698 30200 11704 30252
rect 11756 30240 11762 30252
rect 11756 30212 11801 30240
rect 11756 30200 11762 30212
rect 11882 30200 11888 30252
rect 11940 30200 11946 30252
rect 12158 30249 12164 30252
rect 11977 30243 12035 30249
rect 11977 30209 11989 30243
rect 12023 30209 12035 30243
rect 11977 30203 12035 30209
rect 12115 30243 12164 30249
rect 12115 30209 12127 30243
rect 12161 30209 12164 30243
rect 12115 30203 12164 30209
rect 6733 30175 6791 30181
rect 6733 30172 6745 30175
rect 4571 30144 6040 30172
rect 6564 30144 6745 30172
rect 4571 30141 4583 30144
rect 4525 30135 4583 30141
rect 6012 30104 6040 30144
rect 6733 30141 6745 30144
rect 6779 30172 6791 30175
rect 11992 30172 12020 30203
rect 12158 30200 12164 30203
rect 12216 30200 12222 30252
rect 12342 30200 12348 30252
rect 12400 30240 12406 30252
rect 13722 30240 13728 30252
rect 12400 30212 13728 30240
rect 12400 30200 12406 30212
rect 13722 30200 13728 30212
rect 13780 30200 13786 30252
rect 15194 30200 15200 30252
rect 15252 30240 15258 30252
rect 16114 30240 16120 30252
rect 15252 30212 16120 30240
rect 15252 30200 15258 30212
rect 16114 30200 16120 30212
rect 16172 30200 16178 30252
rect 16482 30200 16488 30252
rect 16540 30240 16546 30252
rect 17681 30243 17739 30249
rect 17681 30240 17693 30243
rect 16540 30212 17693 30240
rect 16540 30200 16546 30212
rect 17681 30209 17693 30212
rect 17727 30209 17739 30243
rect 18417 30243 18475 30249
rect 18417 30240 18429 30243
rect 17681 30203 17739 30209
rect 17880 30212 18429 30240
rect 15286 30172 15292 30184
rect 6779 30144 15292 30172
rect 6779 30141 6791 30144
rect 6733 30135 6791 30141
rect 15286 30132 15292 30144
rect 15344 30172 15350 30184
rect 16666 30172 16672 30184
rect 15344 30144 16672 30172
rect 15344 30132 15350 30144
rect 16666 30132 16672 30144
rect 16724 30132 16730 30184
rect 16758 30132 16764 30184
rect 16816 30172 16822 30184
rect 16942 30172 16948 30184
rect 16816 30144 16948 30172
rect 16816 30132 16822 30144
rect 16942 30132 16948 30144
rect 17000 30132 17006 30184
rect 17218 30132 17224 30184
rect 17276 30172 17282 30184
rect 17773 30175 17831 30181
rect 17773 30172 17785 30175
rect 17276 30144 17785 30172
rect 17276 30132 17282 30144
rect 17773 30141 17785 30144
rect 17819 30141 17831 30175
rect 17773 30135 17831 30141
rect 7469 30107 7527 30113
rect 7469 30104 7481 30107
rect 6012 30076 7481 30104
rect 7469 30073 7481 30076
rect 7515 30073 7527 30107
rect 9490 30104 9496 30116
rect 7469 30067 7527 30073
rect 7576 30076 9496 30104
rect 5258 29996 5264 30048
rect 5316 30036 5322 30048
rect 5718 30036 5724 30048
rect 5316 30008 5724 30036
rect 5316 29996 5322 30008
rect 5718 29996 5724 30008
rect 5776 29996 5782 30048
rect 6822 29996 6828 30048
rect 6880 30036 6886 30048
rect 7576 30036 7604 30076
rect 9490 30064 9496 30076
rect 9548 30064 9554 30116
rect 10686 30064 10692 30116
rect 10744 30104 10750 30116
rect 10744 30076 12434 30104
rect 10744 30064 10750 30076
rect 6880 30008 7604 30036
rect 6880 29996 6886 30008
rect 7926 29996 7932 30048
rect 7984 30036 7990 30048
rect 8665 30039 8723 30045
rect 8665 30036 8677 30039
rect 7984 30008 8677 30036
rect 7984 29996 7990 30008
rect 8665 30005 8677 30008
rect 8711 30036 8723 30039
rect 9398 30036 9404 30048
rect 8711 30008 9404 30036
rect 8711 30005 8723 30008
rect 8665 29999 8723 30005
rect 9398 29996 9404 30008
rect 9456 29996 9462 30048
rect 12250 29996 12256 30048
rect 12308 29996 12314 30048
rect 12406 30036 12434 30076
rect 14550 30064 14556 30116
rect 14608 30104 14614 30116
rect 15838 30104 15844 30116
rect 14608 30076 15844 30104
rect 14608 30064 14614 30076
rect 15838 30064 15844 30076
rect 15896 30064 15902 30116
rect 16684 30104 16712 30132
rect 17880 30104 17908 30212
rect 18417 30209 18429 30212
rect 18463 30209 18475 30243
rect 18417 30203 18475 30209
rect 18506 30200 18512 30252
rect 18564 30200 18570 30252
rect 18598 30200 18604 30252
rect 18656 30200 18662 30252
rect 18785 30243 18843 30249
rect 18785 30209 18797 30243
rect 18831 30209 18843 30243
rect 18785 30203 18843 30209
rect 18322 30132 18328 30184
rect 18380 30172 18386 30184
rect 18690 30172 18696 30184
rect 18380 30144 18696 30172
rect 18380 30132 18386 30144
rect 18690 30132 18696 30144
rect 18748 30172 18754 30184
rect 18800 30172 18828 30203
rect 18966 30200 18972 30252
rect 19024 30200 19030 30252
rect 19058 30200 19064 30252
rect 19116 30240 19122 30252
rect 19904 30240 19932 30271
rect 19978 30268 19984 30280
rect 20036 30268 20042 30320
rect 20088 30317 20116 30348
rect 20257 30345 20269 30379
rect 20303 30376 20315 30379
rect 20346 30376 20352 30388
rect 20303 30348 20352 30376
rect 20303 30345 20315 30348
rect 20257 30339 20315 30345
rect 20346 30336 20352 30348
rect 20404 30336 20410 30388
rect 21082 30336 21088 30388
rect 21140 30376 21146 30388
rect 23842 30376 23848 30388
rect 21140 30348 23848 30376
rect 21140 30336 21146 30348
rect 23842 30336 23848 30348
rect 23900 30336 23906 30388
rect 24688 30348 27108 30376
rect 24688 30320 24716 30348
rect 20073 30311 20131 30317
rect 20073 30277 20085 30311
rect 20119 30277 20131 30311
rect 20441 30311 20499 30317
rect 20441 30308 20453 30311
rect 20073 30271 20131 30277
rect 20272 30280 20453 30308
rect 19116 30212 19932 30240
rect 20272 30240 20300 30280
rect 20441 30277 20453 30280
rect 20487 30277 20499 30311
rect 20441 30271 20499 30277
rect 20622 30268 20628 30320
rect 20680 30308 20686 30320
rect 21174 30308 21180 30320
rect 20680 30280 21180 30308
rect 20680 30268 20686 30280
rect 21174 30268 21180 30280
rect 21232 30268 21238 30320
rect 22646 30268 22652 30320
rect 22704 30308 22710 30320
rect 23198 30308 23204 30320
rect 22704 30280 23204 30308
rect 22704 30268 22710 30280
rect 23198 30268 23204 30280
rect 23256 30268 23262 30320
rect 23382 30268 23388 30320
rect 23440 30268 23446 30320
rect 24670 30268 24676 30320
rect 24728 30268 24734 30320
rect 26602 30308 26608 30320
rect 25700 30280 26608 30308
rect 22002 30240 22008 30252
rect 20272 30212 22008 30240
rect 19116 30200 19122 30212
rect 18748 30144 18828 30172
rect 18984 30172 19012 30200
rect 20272 30172 20300 30212
rect 22002 30200 22008 30212
rect 22060 30200 22066 30252
rect 22922 30200 22928 30252
rect 22980 30240 22986 30252
rect 23106 30240 23112 30252
rect 22980 30212 23112 30240
rect 22980 30200 22986 30212
rect 23106 30200 23112 30212
rect 23164 30200 23170 30252
rect 25700 30249 25728 30280
rect 26602 30268 26608 30280
rect 26660 30268 26666 30320
rect 25685 30243 25743 30249
rect 25685 30240 25697 30243
rect 24688 30212 25697 30240
rect 24688 30172 24716 30212
rect 25685 30209 25697 30212
rect 25731 30209 25743 30243
rect 25685 30203 25743 30209
rect 25774 30200 25780 30252
rect 25832 30240 25838 30252
rect 25869 30243 25927 30249
rect 25869 30240 25881 30243
rect 25832 30212 25881 30240
rect 25832 30200 25838 30212
rect 25869 30209 25881 30212
rect 25915 30209 25927 30243
rect 25869 30203 25927 30209
rect 25958 30200 25964 30252
rect 26016 30200 26022 30252
rect 26053 30243 26111 30249
rect 26053 30209 26065 30243
rect 26099 30240 26111 30243
rect 26142 30240 26148 30252
rect 26099 30212 26148 30240
rect 26099 30209 26111 30212
rect 26053 30203 26111 30209
rect 26142 30200 26148 30212
rect 26200 30200 26206 30252
rect 26234 30200 26240 30252
rect 26292 30240 26298 30252
rect 26510 30240 26516 30252
rect 26292 30212 26516 30240
rect 26292 30200 26298 30212
rect 26510 30200 26516 30212
rect 26568 30200 26574 30252
rect 27080 30240 27108 30348
rect 29086 30336 29092 30388
rect 29144 30336 29150 30388
rect 32950 30376 32956 30388
rect 31726 30348 32956 30376
rect 27798 30268 27804 30320
rect 27856 30308 27862 30320
rect 30650 30308 30656 30320
rect 27856 30280 30656 30308
rect 27856 30268 27862 30280
rect 30650 30268 30656 30280
rect 30708 30308 30714 30320
rect 31018 30308 31024 30320
rect 30708 30280 31024 30308
rect 30708 30268 30714 30280
rect 31018 30268 31024 30280
rect 31076 30268 31082 30320
rect 29822 30240 29828 30252
rect 27080 30212 29828 30240
rect 29822 30200 29828 30212
rect 29880 30200 29886 30252
rect 30377 30243 30435 30249
rect 30377 30209 30389 30243
rect 30423 30240 30435 30243
rect 31294 30240 31300 30252
rect 30423 30212 31300 30240
rect 30423 30209 30435 30212
rect 30377 30203 30435 30209
rect 31294 30200 31300 30212
rect 31352 30200 31358 30252
rect 18984 30144 20300 30172
rect 20364 30144 24716 30172
rect 25133 30175 25191 30181
rect 18748 30132 18754 30144
rect 20364 30116 20392 30144
rect 25133 30141 25145 30175
rect 25179 30172 25191 30175
rect 27338 30172 27344 30184
rect 25179 30144 27344 30172
rect 25179 30141 25191 30144
rect 25133 30135 25191 30141
rect 27338 30132 27344 30144
rect 27396 30132 27402 30184
rect 30834 30132 30840 30184
rect 30892 30172 30898 30184
rect 31726 30172 31754 30348
rect 32950 30336 32956 30348
rect 33008 30376 33014 30388
rect 33008 30348 36032 30376
rect 33008 30336 33014 30348
rect 36004 30320 36032 30348
rect 33042 30308 33048 30320
rect 32416 30280 33048 30308
rect 32030 30200 32036 30252
rect 32088 30240 32094 30252
rect 32125 30243 32183 30249
rect 32125 30240 32137 30243
rect 32088 30212 32137 30240
rect 32088 30200 32094 30212
rect 32125 30209 32137 30212
rect 32171 30209 32183 30243
rect 32125 30203 32183 30209
rect 32306 30200 32312 30252
rect 32364 30200 32370 30252
rect 32416 30249 32444 30280
rect 33042 30268 33048 30280
rect 33100 30308 33106 30320
rect 33226 30308 33232 30320
rect 33100 30280 33232 30308
rect 33100 30268 33106 30280
rect 33226 30268 33232 30280
rect 33284 30268 33290 30320
rect 35986 30268 35992 30320
rect 36044 30268 36050 30320
rect 32401 30243 32459 30249
rect 32401 30209 32413 30243
rect 32447 30209 32459 30243
rect 32401 30203 32459 30209
rect 32490 30200 32496 30252
rect 32548 30200 32554 30252
rect 30892 30144 31754 30172
rect 30892 30132 30898 30144
rect 16684 30076 17908 30104
rect 18049 30107 18107 30113
rect 18049 30073 18061 30107
rect 18095 30104 18107 30107
rect 18095 30076 18460 30104
rect 18095 30073 18107 30076
rect 18049 30067 18107 30073
rect 17402 30036 17408 30048
rect 12406 30008 17408 30036
rect 17402 29996 17408 30008
rect 17460 29996 17466 30048
rect 17862 29996 17868 30048
rect 17920 29996 17926 30048
rect 18141 30039 18199 30045
rect 18141 30005 18153 30039
rect 18187 30036 18199 30039
rect 18322 30036 18328 30048
rect 18187 30008 18328 30036
rect 18187 30005 18199 30008
rect 18141 29999 18199 30005
rect 18322 29996 18328 30008
rect 18380 29996 18386 30048
rect 18432 30036 18460 30076
rect 20346 30064 20352 30116
rect 20404 30064 20410 30116
rect 21542 30104 21548 30116
rect 20640 30076 21548 30104
rect 18690 30036 18696 30048
rect 18432 30008 18696 30036
rect 18690 29996 18696 30008
rect 18748 29996 18754 30048
rect 19886 29996 19892 30048
rect 19944 30036 19950 30048
rect 20073 30039 20131 30045
rect 20073 30036 20085 30039
rect 19944 30008 20085 30036
rect 19944 29996 19950 30008
rect 20073 30005 20085 30008
rect 20119 30036 20131 30039
rect 20438 30036 20444 30048
rect 20119 30008 20444 30036
rect 20119 30005 20131 30008
rect 20073 29999 20131 30005
rect 20438 29996 20444 30008
rect 20496 29996 20502 30048
rect 20530 29996 20536 30048
rect 20588 30036 20594 30048
rect 20640 30045 20668 30076
rect 21542 30064 21548 30076
rect 21600 30064 21606 30116
rect 22278 30064 22284 30116
rect 22336 30104 22342 30116
rect 26050 30104 26056 30116
rect 22336 30076 26056 30104
rect 22336 30064 22342 30076
rect 26050 30064 26056 30076
rect 26108 30064 26114 30116
rect 26602 30064 26608 30116
rect 26660 30104 26666 30116
rect 27798 30104 27804 30116
rect 26660 30076 27804 30104
rect 26660 30064 26666 30076
rect 27798 30064 27804 30076
rect 27856 30064 27862 30116
rect 27982 30064 27988 30116
rect 28040 30104 28046 30116
rect 33318 30104 33324 30116
rect 28040 30076 33324 30104
rect 28040 30064 28046 30076
rect 33318 30064 33324 30076
rect 33376 30064 33382 30116
rect 20625 30039 20683 30045
rect 20625 30036 20637 30039
rect 20588 30008 20637 30036
rect 20588 29996 20594 30008
rect 20625 30005 20637 30008
rect 20671 30005 20683 30039
rect 20625 29999 20683 30005
rect 20806 29996 20812 30048
rect 20864 30036 20870 30048
rect 23934 30036 23940 30048
rect 20864 30008 23940 30036
rect 20864 29996 20870 30008
rect 23934 29996 23940 30008
rect 23992 29996 23998 30048
rect 25314 29996 25320 30048
rect 25372 30036 25378 30048
rect 25774 30036 25780 30048
rect 25372 30008 25780 30036
rect 25372 29996 25378 30008
rect 25774 29996 25780 30008
rect 25832 29996 25838 30048
rect 26237 30039 26295 30045
rect 26237 30005 26249 30039
rect 26283 30036 26295 30039
rect 26694 30036 26700 30048
rect 26283 30008 26700 30036
rect 26283 30005 26295 30008
rect 26237 29999 26295 30005
rect 26694 29996 26700 30008
rect 26752 29996 26758 30048
rect 29914 29996 29920 30048
rect 29972 30036 29978 30048
rect 30558 30036 30564 30048
rect 29972 30008 30564 30036
rect 29972 29996 29978 30008
rect 30558 29996 30564 30008
rect 30616 29996 30622 30048
rect 32769 30039 32827 30045
rect 32769 30005 32781 30039
rect 32815 30036 32827 30039
rect 32950 30036 32956 30048
rect 32815 30008 32956 30036
rect 32815 30005 32827 30008
rect 32769 29999 32827 30005
rect 32950 29996 32956 30008
rect 33008 29996 33014 30048
rect 1104 29946 38272 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38272 29946
rect 1104 29872 38272 29894
rect 10686 29792 10692 29844
rect 10744 29792 10750 29844
rect 12250 29792 12256 29844
rect 12308 29832 12314 29844
rect 12529 29835 12587 29841
rect 12308 29804 12434 29832
rect 12308 29792 12314 29804
rect 6914 29764 6920 29776
rect 4172 29736 6920 29764
rect 3970 29588 3976 29640
rect 4028 29628 4034 29640
rect 4172 29637 4200 29736
rect 6914 29724 6920 29736
rect 6972 29724 6978 29776
rect 8481 29767 8539 29773
rect 8481 29733 8493 29767
rect 8527 29733 8539 29767
rect 8481 29727 8539 29733
rect 6089 29699 6147 29705
rect 6089 29665 6101 29699
rect 6135 29696 6147 29699
rect 6822 29696 6828 29708
rect 6135 29668 6828 29696
rect 6135 29665 6147 29668
rect 6089 29659 6147 29665
rect 6822 29656 6828 29668
rect 6880 29656 6886 29708
rect 8496 29696 8524 29727
rect 9217 29699 9275 29705
rect 9217 29696 9229 29699
rect 8496 29668 9229 29696
rect 9217 29665 9229 29668
rect 9263 29665 9275 29699
rect 12406 29696 12434 29804
rect 12529 29801 12541 29835
rect 12575 29832 12587 29835
rect 12618 29832 12624 29844
rect 12575 29804 12624 29832
rect 12575 29801 12587 29804
rect 12529 29795 12587 29801
rect 12618 29792 12624 29804
rect 12676 29792 12682 29844
rect 15749 29835 15807 29841
rect 15749 29832 15761 29835
rect 14384 29804 15761 29832
rect 14384 29773 14412 29804
rect 15749 29801 15761 29804
rect 15795 29801 15807 29835
rect 15749 29795 15807 29801
rect 16574 29792 16580 29844
rect 16632 29832 16638 29844
rect 16669 29835 16727 29841
rect 16669 29832 16681 29835
rect 16632 29804 16681 29832
rect 16632 29792 16638 29804
rect 16669 29801 16681 29804
rect 16715 29801 16727 29835
rect 16669 29795 16727 29801
rect 17402 29792 17408 29844
rect 17460 29832 17466 29844
rect 17460 29804 19196 29832
rect 17460 29792 17466 29804
rect 13725 29767 13783 29773
rect 13725 29733 13737 29767
rect 13771 29764 13783 29767
rect 14093 29767 14151 29773
rect 14093 29764 14105 29767
rect 13771 29736 14105 29764
rect 13771 29733 13783 29736
rect 13725 29727 13783 29733
rect 14093 29733 14105 29736
rect 14139 29733 14151 29767
rect 14093 29727 14151 29733
rect 14369 29767 14427 29773
rect 14369 29733 14381 29767
rect 14415 29733 14427 29767
rect 15105 29767 15163 29773
rect 15105 29764 15117 29767
rect 14369 29727 14427 29733
rect 14476 29736 15117 29764
rect 14476 29705 14504 29736
rect 15105 29733 15117 29736
rect 15151 29733 15163 29767
rect 15105 29727 15163 29733
rect 15286 29724 15292 29776
rect 15344 29724 15350 29776
rect 18322 29724 18328 29776
rect 18380 29724 18386 29776
rect 18690 29724 18696 29776
rect 18748 29724 18754 29776
rect 18874 29724 18880 29776
rect 18932 29724 18938 29776
rect 19168 29764 19196 29804
rect 19794 29792 19800 29844
rect 19852 29832 19858 29844
rect 20070 29832 20076 29844
rect 19852 29804 20076 29832
rect 19852 29792 19858 29804
rect 20070 29792 20076 29804
rect 20128 29792 20134 29844
rect 20714 29792 20720 29844
rect 20772 29832 20778 29844
rect 21266 29832 21272 29844
rect 20772 29804 21272 29832
rect 20772 29792 20778 29804
rect 21266 29792 21272 29804
rect 21324 29792 21330 29844
rect 22002 29792 22008 29844
rect 22060 29832 22066 29844
rect 24118 29832 24124 29844
rect 22060 29804 24124 29832
rect 22060 29792 22066 29804
rect 24118 29792 24124 29804
rect 24176 29832 24182 29844
rect 24394 29832 24400 29844
rect 24176 29804 24400 29832
rect 24176 29792 24182 29804
rect 24394 29792 24400 29804
rect 24452 29832 24458 29844
rect 24581 29835 24639 29841
rect 24581 29832 24593 29835
rect 24452 29804 24593 29832
rect 24452 29792 24458 29804
rect 24581 29801 24593 29804
rect 24627 29801 24639 29835
rect 24581 29795 24639 29801
rect 25792 29804 31754 29832
rect 20622 29764 20628 29776
rect 19168 29736 20628 29764
rect 20622 29724 20628 29736
rect 20680 29764 20686 29776
rect 23842 29764 23848 29776
rect 20680 29736 21680 29764
rect 20680 29724 20686 29736
rect 14461 29699 14519 29705
rect 12406 29668 13492 29696
rect 9217 29659 9275 29665
rect 4157 29631 4215 29637
rect 4157 29628 4169 29631
rect 4028 29600 4169 29628
rect 4028 29588 4034 29600
rect 4157 29597 4169 29600
rect 4203 29597 4215 29631
rect 4157 29591 4215 29597
rect 5905 29631 5963 29637
rect 5905 29597 5917 29631
rect 5951 29628 5963 29631
rect 5951 29600 6132 29628
rect 5951 29597 5963 29600
rect 5905 29591 5963 29597
rect 6104 29572 6132 29600
rect 8294 29588 8300 29640
rect 8352 29588 8358 29640
rect 8573 29631 8631 29637
rect 8573 29597 8585 29631
rect 8619 29597 8631 29631
rect 8573 29591 8631 29597
rect 8665 29631 8723 29637
rect 8665 29597 8677 29631
rect 8711 29628 8723 29631
rect 8941 29631 8999 29637
rect 8941 29628 8953 29631
rect 8711 29600 8953 29628
rect 8711 29597 8723 29600
rect 8665 29591 8723 29597
rect 8941 29597 8953 29600
rect 8987 29597 8999 29631
rect 8941 29591 8999 29597
rect 5813 29563 5871 29569
rect 5813 29529 5825 29563
rect 5859 29529 5871 29563
rect 5813 29523 5871 29529
rect 4062 29452 4068 29504
rect 4120 29452 4126 29504
rect 5442 29452 5448 29504
rect 5500 29452 5506 29504
rect 5828 29492 5856 29523
rect 6086 29520 6092 29572
rect 6144 29560 6150 29572
rect 8386 29560 8392 29572
rect 6144 29532 8392 29560
rect 6144 29520 6150 29532
rect 8386 29520 8392 29532
rect 8444 29520 8450 29572
rect 6822 29492 6828 29504
rect 5828 29464 6828 29492
rect 6822 29452 6828 29464
rect 6880 29452 6886 29504
rect 8588 29492 8616 29591
rect 12710 29588 12716 29640
rect 12768 29588 12774 29640
rect 13464 29637 13492 29668
rect 14461 29665 14473 29699
rect 14507 29665 14519 29699
rect 15304 29696 15332 29724
rect 18046 29696 18052 29708
rect 15304 29668 15424 29696
rect 14461 29659 14519 29665
rect 12897 29631 12955 29637
rect 12897 29597 12909 29631
rect 12943 29597 12955 29631
rect 12897 29591 12955 29597
rect 13449 29631 13507 29637
rect 13449 29597 13461 29631
rect 13495 29597 13507 29631
rect 13449 29591 13507 29597
rect 9674 29520 9680 29572
rect 9732 29520 9738 29572
rect 12912 29560 12940 29591
rect 13538 29588 13544 29640
rect 13596 29588 13602 29640
rect 13817 29631 13875 29637
rect 13817 29597 13829 29631
rect 13863 29628 13875 29631
rect 13906 29628 13912 29640
rect 13863 29600 13912 29628
rect 13863 29597 13875 29600
rect 13817 29591 13875 29597
rect 13906 29588 13912 29600
rect 13964 29588 13970 29640
rect 14090 29588 14096 29640
rect 14148 29628 14154 29640
rect 14277 29631 14335 29637
rect 14277 29628 14289 29631
rect 14148 29600 14289 29628
rect 14148 29588 14154 29600
rect 14277 29597 14289 29600
rect 14323 29597 14335 29631
rect 14277 29591 14335 29597
rect 14553 29631 14611 29637
rect 14553 29597 14565 29631
rect 14599 29597 14611 29631
rect 14553 29591 14611 29597
rect 14737 29631 14795 29637
rect 14737 29597 14749 29631
rect 14783 29628 14795 29631
rect 14783 29600 15056 29628
rect 14783 29597 14795 29600
rect 14737 29591 14795 29597
rect 14568 29560 14596 29591
rect 15028 29572 15056 29600
rect 15102 29588 15108 29640
rect 15160 29628 15166 29640
rect 15396 29637 15424 29668
rect 15948 29668 18052 29696
rect 15289 29631 15347 29637
rect 15289 29628 15301 29631
rect 15160 29600 15301 29628
rect 15160 29588 15166 29600
rect 15289 29597 15301 29600
rect 15335 29597 15347 29631
rect 15289 29591 15347 29597
rect 15381 29631 15439 29637
rect 15381 29597 15393 29631
rect 15427 29597 15439 29631
rect 15381 29591 15439 29597
rect 15470 29588 15476 29640
rect 15528 29588 15534 29640
rect 15654 29588 15660 29640
rect 15712 29588 15718 29640
rect 15838 29588 15844 29640
rect 15896 29628 15902 29640
rect 15948 29637 15976 29668
rect 18046 29656 18052 29668
rect 18104 29656 18110 29708
rect 15933 29631 15991 29637
rect 15933 29628 15945 29631
rect 15896 29600 15945 29628
rect 15896 29588 15902 29600
rect 15933 29597 15945 29600
rect 15979 29597 15991 29631
rect 15933 29591 15991 29597
rect 16114 29588 16120 29640
rect 16172 29588 16178 29640
rect 16301 29631 16359 29637
rect 16301 29597 16313 29631
rect 16347 29628 16359 29631
rect 16347 29600 17264 29628
rect 16347 29597 16359 29600
rect 16301 29591 16359 29597
rect 12912 29532 14596 29560
rect 9030 29492 9036 29504
rect 8588 29464 9036 29492
rect 9030 29452 9036 29464
rect 9088 29492 9094 29504
rect 9950 29492 9956 29504
rect 9088 29464 9956 29492
rect 9088 29452 9094 29464
rect 9950 29452 9956 29464
rect 10008 29452 10014 29504
rect 13262 29452 13268 29504
rect 13320 29452 13326 29504
rect 14568 29492 14596 29532
rect 15010 29520 15016 29572
rect 15068 29520 15074 29572
rect 16022 29520 16028 29572
rect 16080 29520 16086 29572
rect 16132 29560 16160 29588
rect 16390 29560 16396 29572
rect 16132 29532 16396 29560
rect 16390 29520 16396 29532
rect 16448 29520 16454 29572
rect 17236 29569 17264 29600
rect 18138 29588 18144 29640
rect 18196 29628 18202 29640
rect 18340 29637 18368 29724
rect 18708 29696 18736 29724
rect 21652 29708 21680 29736
rect 23252 29736 23848 29764
rect 18616 29668 18736 29696
rect 18233 29631 18291 29637
rect 18233 29628 18245 29631
rect 18196 29600 18245 29628
rect 18196 29588 18202 29600
rect 18233 29597 18245 29600
rect 18279 29597 18291 29631
rect 18233 29591 18291 29597
rect 18325 29631 18383 29637
rect 18325 29597 18337 29631
rect 18371 29597 18383 29631
rect 18325 29591 18383 29597
rect 18506 29588 18512 29640
rect 18564 29588 18570 29640
rect 18616 29637 18644 29668
rect 18966 29656 18972 29708
rect 19024 29696 19030 29708
rect 19702 29696 19708 29708
rect 19024 29668 19708 29696
rect 19024 29656 19030 29668
rect 19702 29656 19708 29668
rect 19760 29656 19766 29708
rect 19886 29656 19892 29708
rect 19944 29696 19950 29708
rect 19944 29668 20668 29696
rect 19944 29656 19950 29668
rect 18601 29631 18659 29637
rect 18601 29597 18613 29631
rect 18647 29597 18659 29631
rect 18601 29591 18659 29597
rect 18690 29588 18696 29640
rect 18748 29588 18754 29640
rect 19150 29588 19156 29640
rect 19208 29628 19214 29640
rect 20530 29628 20536 29640
rect 19208 29600 20536 29628
rect 19208 29588 19214 29600
rect 20530 29588 20536 29600
rect 20588 29588 20594 29640
rect 20640 29628 20668 29668
rect 21634 29656 21640 29708
rect 21692 29656 21698 29708
rect 22756 29668 23152 29696
rect 22756 29640 22784 29668
rect 20901 29631 20959 29637
rect 20640 29625 20760 29628
rect 20901 29625 20913 29631
rect 20640 29600 20913 29625
rect 20732 29597 20913 29600
rect 20947 29597 20959 29631
rect 20901 29591 20959 29597
rect 20993 29631 21051 29637
rect 20993 29597 21005 29631
rect 21039 29628 21051 29631
rect 21266 29628 21272 29640
rect 21039 29600 21272 29628
rect 21039 29597 21051 29600
rect 20993 29591 21051 29597
rect 21266 29588 21272 29600
rect 21324 29588 21330 29640
rect 21450 29588 21456 29640
rect 21508 29628 21514 29640
rect 21508 29600 22416 29628
rect 21508 29588 21514 29600
rect 17221 29563 17279 29569
rect 17221 29529 17233 29563
rect 17267 29529 17279 29563
rect 22278 29560 22284 29572
rect 17221 29523 17279 29529
rect 19260 29532 22284 29560
rect 16758 29492 16764 29504
rect 14568 29464 16764 29492
rect 16758 29452 16764 29464
rect 16816 29452 16822 29504
rect 16850 29452 16856 29504
rect 16908 29452 16914 29504
rect 16942 29452 16948 29504
rect 17000 29452 17006 29504
rect 17034 29452 17040 29504
rect 17092 29452 17098 29504
rect 17236 29492 17264 29523
rect 19260 29492 19288 29532
rect 22278 29520 22284 29532
rect 22336 29520 22342 29572
rect 22388 29560 22416 29600
rect 22738 29588 22744 29640
rect 22796 29588 22802 29640
rect 22922 29637 22928 29640
rect 22920 29628 22928 29637
rect 22883 29600 22928 29628
rect 22920 29591 22928 29600
rect 22922 29588 22928 29591
rect 22980 29588 22986 29640
rect 23124 29637 23152 29668
rect 23252 29640 23280 29736
rect 23842 29724 23848 29736
rect 23900 29724 23906 29776
rect 25130 29764 25136 29776
rect 24044 29736 25136 29764
rect 23474 29656 23480 29708
rect 23532 29696 23538 29708
rect 23532 29668 23796 29696
rect 23532 29656 23538 29668
rect 23768 29640 23796 29668
rect 23109 29631 23167 29637
rect 23109 29597 23121 29631
rect 23155 29597 23167 29631
rect 23109 29591 23167 29597
rect 23198 29588 23204 29640
rect 23256 29637 23280 29640
rect 23256 29631 23295 29637
rect 23283 29597 23295 29631
rect 23256 29591 23295 29597
rect 23256 29588 23262 29591
rect 23382 29588 23388 29640
rect 23440 29588 23446 29640
rect 23750 29588 23756 29640
rect 23808 29588 23814 29640
rect 24044 29637 24072 29736
rect 25130 29724 25136 29736
rect 25188 29724 25194 29776
rect 24578 29656 24584 29708
rect 24636 29656 24642 29708
rect 24670 29656 24676 29708
rect 24728 29656 24734 29708
rect 24029 29631 24087 29637
rect 24029 29597 24041 29631
rect 24075 29597 24087 29631
rect 24029 29591 24087 29597
rect 24302 29588 24308 29640
rect 24360 29628 24366 29640
rect 24596 29628 24624 29656
rect 24765 29631 24823 29637
rect 24765 29628 24777 29631
rect 24360 29600 24777 29628
rect 24360 29588 24366 29600
rect 24765 29597 24777 29600
rect 24811 29597 24823 29631
rect 24765 29591 24823 29597
rect 23017 29563 23075 29569
rect 23017 29560 23029 29563
rect 22388 29532 23029 29560
rect 23017 29529 23029 29532
rect 23063 29529 23075 29563
rect 24780 29560 24808 29591
rect 24946 29588 24952 29640
rect 25004 29628 25010 29640
rect 25792 29637 25820 29804
rect 26050 29724 26056 29776
rect 26108 29764 26114 29776
rect 26108 29736 26556 29764
rect 26108 29724 26114 29736
rect 26237 29699 26295 29705
rect 26237 29696 26249 29699
rect 25976 29668 26249 29696
rect 25976 29637 26004 29668
rect 26237 29665 26249 29668
rect 26283 29665 26295 29699
rect 26237 29659 26295 29665
rect 25777 29631 25835 29637
rect 25777 29628 25789 29631
rect 25004 29600 25789 29628
rect 25004 29588 25010 29600
rect 25777 29597 25789 29600
rect 25823 29597 25835 29631
rect 25777 29591 25835 29597
rect 25869 29631 25927 29637
rect 25869 29597 25881 29631
rect 25915 29597 25927 29631
rect 25869 29591 25927 29597
rect 25961 29631 26019 29637
rect 25961 29597 25973 29631
rect 26007 29597 26019 29631
rect 25961 29591 26019 29597
rect 25884 29560 25912 29591
rect 26050 29588 26056 29640
rect 26108 29628 26114 29640
rect 26145 29631 26203 29637
rect 26145 29628 26157 29631
rect 26108 29600 26157 29628
rect 26108 29588 26114 29600
rect 26145 29597 26157 29600
rect 26191 29628 26203 29631
rect 26326 29628 26332 29640
rect 26191 29600 26332 29628
rect 26191 29597 26203 29600
rect 26145 29591 26203 29597
rect 26326 29588 26332 29600
rect 26384 29588 26390 29640
rect 26418 29588 26424 29640
rect 26476 29588 26482 29640
rect 26528 29637 26556 29736
rect 26694 29724 26700 29776
rect 26752 29724 26758 29776
rect 27338 29724 27344 29776
rect 27396 29764 27402 29776
rect 28718 29764 28724 29776
rect 27396 29736 28724 29764
rect 27396 29724 27402 29736
rect 28718 29724 28724 29736
rect 28776 29724 28782 29776
rect 29270 29724 29276 29776
rect 29328 29764 29334 29776
rect 30374 29764 30380 29776
rect 29328 29736 30380 29764
rect 29328 29724 29334 29736
rect 30374 29724 30380 29736
rect 30432 29764 30438 29776
rect 30432 29736 30512 29764
rect 30432 29724 30438 29736
rect 26712 29637 26740 29724
rect 27356 29696 27384 29724
rect 27356 29668 27476 29696
rect 26513 29631 26571 29637
rect 26513 29597 26525 29631
rect 26559 29597 26571 29631
rect 26513 29591 26571 29597
rect 26697 29631 26755 29637
rect 26697 29597 26709 29631
rect 26743 29597 26755 29631
rect 26697 29591 26755 29597
rect 24780 29532 25912 29560
rect 26528 29560 26556 29591
rect 26786 29588 26792 29640
rect 26844 29588 26850 29640
rect 27338 29588 27344 29640
rect 27396 29588 27402 29640
rect 27448 29637 27476 29668
rect 27614 29656 27620 29708
rect 27672 29656 27678 29708
rect 28994 29696 29000 29708
rect 27816 29668 29000 29696
rect 27433 29631 27491 29637
rect 27433 29597 27445 29631
rect 27479 29597 27491 29631
rect 27433 29591 27491 29597
rect 26528 29532 26648 29560
rect 23017 29523 23075 29529
rect 17236 29464 19288 29492
rect 20809 29495 20867 29501
rect 20809 29461 20821 29495
rect 20855 29492 20867 29495
rect 20990 29492 20996 29504
rect 20855 29464 20996 29492
rect 20855 29461 20867 29464
rect 20809 29455 20867 29461
rect 20990 29452 20996 29464
rect 21048 29452 21054 29504
rect 21177 29495 21235 29501
rect 21177 29461 21189 29495
rect 21223 29492 21235 29495
rect 21818 29492 21824 29504
rect 21223 29464 21824 29492
rect 21223 29461 21235 29464
rect 21177 29455 21235 29461
rect 21818 29452 21824 29464
rect 21876 29452 21882 29504
rect 22646 29452 22652 29504
rect 22704 29492 22710 29504
rect 22741 29495 22799 29501
rect 22741 29492 22753 29495
rect 22704 29464 22753 29492
rect 22704 29452 22710 29464
rect 22741 29461 22753 29464
rect 22787 29461 22799 29495
rect 23032 29492 23060 29523
rect 23290 29492 23296 29504
rect 23032 29464 23296 29492
rect 22741 29455 22799 29461
rect 23290 29452 23296 29464
rect 23348 29452 23354 29504
rect 23566 29452 23572 29504
rect 23624 29452 23630 29504
rect 23937 29495 23995 29501
rect 23937 29461 23949 29495
rect 23983 29492 23995 29495
rect 24397 29495 24455 29501
rect 24397 29492 24409 29495
rect 23983 29464 24409 29492
rect 23983 29461 23995 29464
rect 23937 29455 23995 29461
rect 24397 29461 24409 29464
rect 24443 29461 24455 29495
rect 24397 29455 24455 29461
rect 25501 29495 25559 29501
rect 25501 29461 25513 29495
rect 25547 29492 25559 29495
rect 25774 29492 25780 29504
rect 25547 29464 25780 29492
rect 25547 29461 25559 29464
rect 25501 29455 25559 29461
rect 25774 29452 25780 29464
rect 25832 29452 25838 29504
rect 25884 29492 25912 29532
rect 26510 29492 26516 29504
rect 25884 29464 26516 29492
rect 26510 29452 26516 29464
rect 26568 29452 26574 29504
rect 26620 29492 26648 29532
rect 27816 29501 27844 29668
rect 28994 29656 29000 29668
rect 29052 29696 29058 29708
rect 29052 29668 30420 29696
rect 29052 29656 29058 29668
rect 28537 29631 28595 29637
rect 28537 29628 28549 29631
rect 28184 29600 28549 29628
rect 27801 29495 27859 29501
rect 27801 29492 27813 29495
rect 26620 29464 27813 29492
rect 27801 29461 27813 29464
rect 27847 29461 27859 29495
rect 27801 29455 27859 29461
rect 27893 29495 27951 29501
rect 27893 29461 27905 29495
rect 27939 29492 27951 29495
rect 27982 29492 27988 29504
rect 27939 29464 27988 29492
rect 27939 29461 27951 29464
rect 27893 29455 27951 29461
rect 27982 29452 27988 29464
rect 28040 29452 28046 29504
rect 28184 29492 28212 29600
rect 28537 29597 28549 29600
rect 28583 29597 28595 29631
rect 28537 29591 28595 29597
rect 28718 29588 28724 29640
rect 28776 29628 28782 29640
rect 29365 29631 29423 29637
rect 29365 29628 29377 29631
rect 28776 29600 29377 29628
rect 28776 29588 28782 29600
rect 29365 29597 29377 29600
rect 29411 29628 29423 29631
rect 29638 29628 29644 29640
rect 29411 29600 29644 29628
rect 29411 29597 29423 29600
rect 29365 29591 29423 29597
rect 29638 29588 29644 29600
rect 29696 29588 29702 29640
rect 29822 29588 29828 29640
rect 29880 29588 29886 29640
rect 29917 29631 29975 29637
rect 29917 29597 29929 29631
rect 29963 29597 29975 29631
rect 29917 29591 29975 29597
rect 28261 29495 28319 29501
rect 28261 29492 28273 29495
rect 28184 29464 28273 29492
rect 28261 29461 28273 29464
rect 28307 29461 28319 29495
rect 28261 29455 28319 29461
rect 28350 29452 28356 29504
rect 28408 29452 28414 29504
rect 29270 29452 29276 29504
rect 29328 29452 29334 29504
rect 29546 29452 29552 29504
rect 29604 29452 29610 29504
rect 29822 29452 29828 29504
rect 29880 29492 29886 29504
rect 29932 29492 29960 29591
rect 30006 29588 30012 29640
rect 30064 29588 30070 29640
rect 30190 29588 30196 29640
rect 30248 29588 30254 29640
rect 30392 29637 30420 29668
rect 30285 29631 30343 29637
rect 30285 29597 30297 29631
rect 30331 29597 30343 29631
rect 30285 29591 30343 29597
rect 30378 29631 30436 29637
rect 30378 29597 30390 29631
rect 30424 29597 30436 29631
rect 30378 29591 30436 29597
rect 30300 29560 30328 29591
rect 30484 29560 30512 29736
rect 31726 29640 31754 29804
rect 34054 29764 34060 29776
rect 33980 29736 34060 29764
rect 33980 29705 34008 29736
rect 34054 29724 34060 29736
rect 34112 29764 34118 29776
rect 34238 29764 34244 29776
rect 34112 29736 34244 29764
rect 34112 29724 34118 29736
rect 34238 29724 34244 29736
rect 34296 29724 34302 29776
rect 33965 29699 34023 29705
rect 33965 29665 33977 29699
rect 34011 29665 34023 29699
rect 36817 29699 36875 29705
rect 36817 29696 36829 29699
rect 33965 29659 34023 29665
rect 34164 29668 36829 29696
rect 30558 29588 30564 29640
rect 30616 29588 30622 29640
rect 30742 29588 30748 29640
rect 30800 29637 30806 29640
rect 30800 29631 30849 29637
rect 30800 29597 30803 29631
rect 30837 29628 30849 29631
rect 31018 29628 31024 29640
rect 30837 29600 31024 29628
rect 30837 29597 30849 29600
rect 30800 29591 30849 29597
rect 30800 29588 30806 29591
rect 31018 29588 31024 29600
rect 31076 29588 31082 29640
rect 31205 29631 31263 29637
rect 31205 29597 31217 29631
rect 31251 29628 31263 29631
rect 31294 29628 31300 29640
rect 31251 29600 31300 29628
rect 31251 29597 31263 29600
rect 31205 29591 31263 29597
rect 31294 29588 31300 29600
rect 31352 29588 31358 29640
rect 31662 29588 31668 29640
rect 31720 29628 31754 29640
rect 34164 29637 34192 29668
rect 36817 29665 36829 29668
rect 36863 29665 36875 29699
rect 36817 29659 36875 29665
rect 34149 29631 34207 29637
rect 34149 29628 34161 29631
rect 31720 29600 34161 29628
rect 31720 29588 31726 29600
rect 34149 29597 34161 29600
rect 34195 29597 34207 29631
rect 34149 29591 34207 29597
rect 34790 29588 34796 29640
rect 34848 29588 34854 29640
rect 30300 29532 30512 29560
rect 30650 29520 30656 29572
rect 30708 29520 30714 29572
rect 31110 29560 31116 29572
rect 30852 29532 31116 29560
rect 30852 29492 30880 29532
rect 31110 29520 31116 29532
rect 31168 29520 31174 29572
rect 32953 29563 33011 29569
rect 32953 29529 32965 29563
rect 32999 29560 33011 29563
rect 34330 29560 34336 29572
rect 32999 29532 34336 29560
rect 32999 29529 33011 29532
rect 32953 29523 33011 29529
rect 34330 29520 34336 29532
rect 34388 29520 34394 29572
rect 34974 29520 34980 29572
rect 35032 29560 35038 29572
rect 35069 29563 35127 29569
rect 35069 29560 35081 29563
rect 35032 29532 35081 29560
rect 35032 29520 35038 29532
rect 35069 29529 35081 29532
rect 35115 29529 35127 29563
rect 35069 29523 35127 29529
rect 29880 29464 30880 29492
rect 29880 29452 29886 29464
rect 30926 29452 30932 29504
rect 30984 29452 30990 29504
rect 33318 29452 33324 29504
rect 33376 29492 33382 29504
rect 34057 29495 34115 29501
rect 34057 29492 34069 29495
rect 33376 29464 34069 29492
rect 33376 29452 33382 29464
rect 34057 29461 34069 29464
rect 34103 29461 34115 29495
rect 34057 29455 34115 29461
rect 34514 29452 34520 29504
rect 34572 29452 34578 29504
rect 35986 29452 35992 29504
rect 36044 29492 36050 29504
rect 36188 29492 36216 29614
rect 36044 29464 36216 29492
rect 36044 29452 36050 29464
rect 1104 29402 38272 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38272 29402
rect 1104 29328 38272 29350
rect 4062 29248 4068 29300
rect 4120 29248 4126 29300
rect 6822 29248 6828 29300
rect 6880 29288 6886 29300
rect 6880 29260 7052 29288
rect 6880 29248 6886 29260
rect 4080 29220 4108 29248
rect 3896 29192 4108 29220
rect 3896 29161 3924 29192
rect 6086 29180 6092 29232
rect 6144 29180 6150 29232
rect 7024 29229 7052 29260
rect 8294 29248 8300 29300
rect 8352 29288 8358 29300
rect 8757 29291 8815 29297
rect 8757 29288 8769 29291
rect 8352 29260 8769 29288
rect 8352 29248 8358 29260
rect 8757 29257 8769 29260
rect 8803 29257 8815 29291
rect 8757 29251 8815 29257
rect 9125 29291 9183 29297
rect 9125 29257 9137 29291
rect 9171 29288 9183 29291
rect 10686 29288 10692 29300
rect 9171 29260 10692 29288
rect 9171 29257 9183 29260
rect 9125 29251 9183 29257
rect 10686 29248 10692 29260
rect 10744 29248 10750 29300
rect 16758 29248 16764 29300
rect 16816 29288 16822 29300
rect 16816 29260 18092 29288
rect 16816 29248 16822 29260
rect 7009 29223 7067 29229
rect 7009 29189 7021 29223
rect 7055 29220 7067 29223
rect 11333 29223 11391 29229
rect 7055 29192 9168 29220
rect 7055 29189 7067 29192
rect 7009 29183 7067 29189
rect 3881 29155 3939 29161
rect 3881 29121 3893 29155
rect 3927 29121 3939 29155
rect 3881 29115 3939 29121
rect 5258 29112 5264 29164
rect 5316 29152 5322 29164
rect 5316 29124 5396 29152
rect 5316 29112 5322 29124
rect 5368 28960 5396 29124
rect 5905 29087 5963 29093
rect 5905 29053 5917 29087
rect 5951 29084 5963 29087
rect 6104 29084 6132 29180
rect 6917 29155 6975 29161
rect 6917 29121 6929 29155
rect 6963 29121 6975 29155
rect 6917 29115 6975 29121
rect 7101 29155 7159 29161
rect 7101 29121 7113 29155
rect 7147 29121 7159 29155
rect 7101 29115 7159 29121
rect 7285 29155 7343 29161
rect 7285 29121 7297 29155
rect 7331 29152 7343 29155
rect 7653 29155 7711 29161
rect 7653 29152 7665 29155
rect 7331 29124 7665 29152
rect 7331 29121 7343 29124
rect 7285 29115 7343 29121
rect 7653 29121 7665 29124
rect 7699 29121 7711 29155
rect 7653 29115 7711 29121
rect 5951 29056 6132 29084
rect 6932 29084 6960 29115
rect 7006 29084 7012 29096
rect 6932 29056 7012 29084
rect 5951 29053 5963 29056
rect 5905 29047 5963 29053
rect 7006 29044 7012 29056
rect 7064 29044 7070 29096
rect 7116 29084 7144 29115
rect 7926 29112 7932 29164
rect 7984 29112 7990 29164
rect 8128 29124 8432 29152
rect 7944 29084 7972 29112
rect 7116 29056 7972 29084
rect 6914 28976 6920 29028
rect 6972 29016 6978 29028
rect 8128 29016 8156 29124
rect 8297 29087 8355 29093
rect 8297 29084 8309 29087
rect 6972 28988 8156 29016
rect 8220 29056 8309 29084
rect 8220 28994 8248 29056
rect 8297 29053 8309 29056
rect 8343 29053 8355 29087
rect 8297 29047 8355 29053
rect 8404 29016 8432 29124
rect 9140 29096 9168 29192
rect 11333 29189 11345 29223
rect 11379 29220 11391 29223
rect 17954 29220 17960 29232
rect 11379 29192 17960 29220
rect 11379 29189 11391 29192
rect 11333 29183 11391 29189
rect 17954 29180 17960 29192
rect 18012 29180 18018 29232
rect 18064 29220 18092 29260
rect 18690 29248 18696 29300
rect 18748 29288 18754 29300
rect 18877 29291 18935 29297
rect 18877 29288 18889 29291
rect 18748 29260 18889 29288
rect 18748 29248 18754 29260
rect 18877 29257 18889 29260
rect 18923 29257 18935 29291
rect 18877 29251 18935 29257
rect 18966 29248 18972 29300
rect 19024 29248 19030 29300
rect 21450 29288 21456 29300
rect 21008 29260 21456 29288
rect 18064 29192 18736 29220
rect 12710 29112 12716 29164
rect 12768 29152 12774 29164
rect 13081 29155 13139 29161
rect 13081 29152 13093 29155
rect 12768 29124 13093 29152
rect 12768 29112 12774 29124
rect 13081 29121 13093 29124
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 13265 29155 13323 29161
rect 13265 29121 13277 29155
rect 13311 29152 13323 29155
rect 16666 29152 16672 29164
rect 13311 29124 16672 29152
rect 13311 29121 13323 29124
rect 13265 29115 13323 29121
rect 16666 29112 16672 29124
rect 16724 29112 16730 29164
rect 16850 29112 16856 29164
rect 16908 29152 16914 29164
rect 17218 29152 17224 29164
rect 16908 29124 17224 29152
rect 16908 29112 16914 29124
rect 17218 29112 17224 29124
rect 17276 29152 17282 29164
rect 17494 29152 17500 29164
rect 17276 29124 17500 29152
rect 17276 29112 17282 29124
rect 17494 29112 17500 29124
rect 17552 29112 17558 29164
rect 17678 29112 17684 29164
rect 17736 29152 17742 29164
rect 18414 29152 18420 29164
rect 17736 29124 18420 29152
rect 17736 29112 17742 29124
rect 18414 29112 18420 29124
rect 18472 29112 18478 29164
rect 18509 29155 18567 29161
rect 18509 29121 18521 29155
rect 18555 29152 18567 29155
rect 18598 29152 18604 29164
rect 18555 29124 18604 29152
rect 18555 29121 18567 29124
rect 18509 29115 18567 29121
rect 18598 29112 18604 29124
rect 18656 29112 18662 29164
rect 18708 29161 18736 29192
rect 18693 29155 18751 29161
rect 18693 29121 18705 29155
rect 18739 29152 18751 29155
rect 18984 29152 19012 29248
rect 20346 29220 20352 29232
rect 18739 29124 19012 29152
rect 19260 29192 20352 29220
rect 18739 29121 18751 29124
rect 18693 29115 18751 29121
rect 9122 29044 9128 29096
rect 9180 29084 9186 29096
rect 9217 29087 9275 29093
rect 9217 29084 9229 29087
rect 9180 29056 9229 29084
rect 9180 29044 9186 29056
rect 9217 29053 9229 29056
rect 9263 29053 9275 29087
rect 9217 29047 9275 29053
rect 9401 29087 9459 29093
rect 9401 29053 9413 29087
rect 9447 29084 9459 29087
rect 10962 29084 10968 29096
rect 9447 29056 10968 29084
rect 9447 29053 9459 29056
rect 9401 29047 9459 29053
rect 10962 29044 10968 29056
rect 11020 29044 11026 29096
rect 16022 29044 16028 29096
rect 16080 29084 16086 29096
rect 19260 29084 19288 29192
rect 20346 29180 20352 29192
rect 20404 29180 20410 29232
rect 20898 29180 20904 29232
rect 20956 29180 20962 29232
rect 19886 29112 19892 29164
rect 19944 29112 19950 29164
rect 20622 29112 20628 29164
rect 20680 29158 20686 29164
rect 21008 29161 21036 29260
rect 21450 29248 21456 29260
rect 21508 29248 21514 29300
rect 21634 29248 21640 29300
rect 21692 29288 21698 29300
rect 21692 29260 23796 29288
rect 21692 29248 21698 29260
rect 22370 29220 22376 29232
rect 21652 29192 22376 29220
rect 21652 29164 21680 29192
rect 20717 29158 20775 29161
rect 20680 29155 20775 29158
rect 20680 29130 20729 29155
rect 20680 29112 20686 29130
rect 20717 29121 20729 29130
rect 20763 29121 20775 29155
rect 20993 29155 21051 29161
rect 20993 29152 21005 29155
rect 20717 29115 20775 29121
rect 20917 29124 21005 29152
rect 16080 29056 19288 29084
rect 19904 29084 19932 29112
rect 20917 29084 20945 29124
rect 20993 29121 21005 29124
rect 21039 29121 21051 29155
rect 20993 29115 21051 29121
rect 21082 29112 21088 29164
rect 21140 29112 21146 29164
rect 21634 29112 21640 29164
rect 21692 29112 21698 29164
rect 21818 29112 21824 29164
rect 21876 29112 21882 29164
rect 22002 29161 22008 29164
rect 21969 29155 22008 29161
rect 21969 29121 21981 29155
rect 21969 29115 22008 29121
rect 22002 29112 22008 29115
rect 22060 29112 22066 29164
rect 22094 29112 22100 29164
rect 22152 29112 22158 29164
rect 22186 29112 22192 29164
rect 22244 29112 22250 29164
rect 22293 29161 22321 29192
rect 22370 29180 22376 29192
rect 22428 29180 22434 29232
rect 23198 29180 23204 29232
rect 23256 29220 23262 29232
rect 23256 29192 23520 29220
rect 23256 29180 23262 29192
rect 22286 29155 22344 29161
rect 22286 29121 22298 29155
rect 22332 29121 22344 29155
rect 22286 29115 22344 29121
rect 22554 29112 22560 29164
rect 22612 29112 22618 29164
rect 22646 29112 22652 29164
rect 22704 29152 22710 29164
rect 22833 29155 22891 29161
rect 22833 29152 22845 29155
rect 22704 29124 22845 29152
rect 22704 29112 22710 29124
rect 22833 29121 22845 29124
rect 22879 29121 22891 29155
rect 22833 29115 22891 29121
rect 23014 29112 23020 29164
rect 23072 29112 23078 29164
rect 23492 29161 23520 29192
rect 23658 29180 23664 29232
rect 23716 29180 23722 29232
rect 23768 29161 23796 29260
rect 23842 29248 23848 29300
rect 23900 29288 23906 29300
rect 26418 29288 26424 29300
rect 23900 29260 25820 29288
rect 23900 29248 23906 29260
rect 23477 29155 23535 29161
rect 23477 29121 23489 29155
rect 23523 29121 23535 29155
rect 23477 29115 23535 29121
rect 23753 29155 23811 29161
rect 23753 29121 23765 29155
rect 23799 29121 23811 29155
rect 23753 29115 23811 29121
rect 23845 29155 23903 29161
rect 23845 29121 23857 29155
rect 23891 29152 23903 29155
rect 23934 29152 23940 29164
rect 23891 29124 23940 29152
rect 23891 29121 23903 29124
rect 23845 29115 23903 29121
rect 23934 29112 23940 29124
rect 23992 29112 23998 29164
rect 25406 29112 25412 29164
rect 25464 29152 25470 29164
rect 25501 29155 25559 29161
rect 25501 29152 25513 29155
rect 25464 29124 25513 29152
rect 25464 29112 25470 29124
rect 25501 29121 25513 29124
rect 25547 29121 25559 29155
rect 25501 29115 25559 29121
rect 19904 29056 20945 29084
rect 16080 29044 16086 29056
rect 9861 29019 9919 29025
rect 9861 29016 9873 29019
rect 6972 28976 6978 28988
rect 8220 28966 8340 28994
rect 8404 28988 9873 29016
rect 9861 28985 9873 28988
rect 9907 28985 9919 29019
rect 9861 28979 9919 28985
rect 12894 28976 12900 29028
rect 12952 28976 12958 29028
rect 13722 28976 13728 29028
rect 13780 29016 13786 29028
rect 13780 28988 20945 29016
rect 13780 28976 13786 28988
rect 4144 28951 4202 28957
rect 4144 28917 4156 28951
rect 4190 28948 4202 28951
rect 4614 28948 4620 28960
rect 4190 28920 4620 28948
rect 4190 28917 4202 28920
rect 4144 28911 4202 28917
rect 4614 28908 4620 28920
rect 4672 28908 4678 28960
rect 5350 28908 5356 28960
rect 5408 28908 5414 28960
rect 6546 28908 6552 28960
rect 6604 28948 6610 28960
rect 6733 28951 6791 28957
rect 6733 28948 6745 28951
rect 6604 28920 6745 28948
rect 6604 28908 6610 28920
rect 6733 28917 6745 28920
rect 6779 28917 6791 28951
rect 8312 28948 8340 28966
rect 8386 28948 8392 28960
rect 8312 28920 8392 28948
rect 6733 28911 6791 28917
rect 8386 28908 8392 28920
rect 8444 28908 8450 28960
rect 8478 28908 8484 28960
rect 8536 28948 8542 28960
rect 18414 28948 18420 28960
rect 8536 28920 18420 28948
rect 8536 28908 8542 28920
rect 18414 28908 18420 28920
rect 18472 28908 18478 28960
rect 18598 28908 18604 28960
rect 18656 28908 18662 28960
rect 19150 28908 19156 28960
rect 19208 28948 19214 28960
rect 19886 28948 19892 28960
rect 19208 28920 19892 28948
rect 19208 28908 19214 28920
rect 19886 28908 19892 28920
rect 19944 28908 19950 28960
rect 20917 28948 20945 28988
rect 21100 28948 21128 29112
rect 22741 29087 22799 29093
rect 22741 29053 22753 29087
rect 22787 29084 22799 29087
rect 22787 29056 23336 29084
rect 22787 29053 22799 29056
rect 22741 29047 22799 29053
rect 22465 29019 22523 29025
rect 21266 28994 21272 29006
rect 21225 28966 21272 28994
rect 21266 28954 21272 28966
rect 21324 28954 21330 29006
rect 22465 28985 22477 29019
rect 22511 29016 22523 29019
rect 22925 29019 22983 29025
rect 22925 29016 22937 29019
rect 22511 28988 22937 29016
rect 22511 28985 22523 28988
rect 22465 28979 22523 28985
rect 22925 28985 22937 28988
rect 22971 28985 22983 29019
rect 23308 29016 23336 29056
rect 23934 29016 23940 29028
rect 23308 28988 23428 29016
rect 22925 28979 22983 28985
rect 20917 28920 21128 28948
rect 21269 28951 21327 28954
rect 21269 28917 21281 28951
rect 21315 28917 21327 28951
rect 21269 28911 21327 28917
rect 23198 28908 23204 28960
rect 23256 28908 23262 28960
rect 23400 28948 23428 28988
rect 23584 28988 23940 29016
rect 23584 28948 23612 28988
rect 23934 28976 23940 28988
rect 23992 28976 23998 29028
rect 25516 29016 25544 29115
rect 25590 29112 25596 29164
rect 25648 29112 25654 29164
rect 25792 29161 25820 29260
rect 25884 29260 26424 29288
rect 25884 29161 25912 29260
rect 26418 29248 26424 29260
rect 26476 29248 26482 29300
rect 26510 29248 26516 29300
rect 26568 29248 26574 29300
rect 27338 29248 27344 29300
rect 27396 29248 27402 29300
rect 28350 29288 28356 29300
rect 27908 29260 28356 29288
rect 26053 29223 26111 29229
rect 26053 29189 26065 29223
rect 26099 29220 26111 29223
rect 26528 29220 26556 29248
rect 27356 29220 27384 29248
rect 26099 29192 26372 29220
rect 26099 29189 26111 29192
rect 26053 29183 26111 29189
rect 25777 29155 25835 29161
rect 25777 29121 25789 29155
rect 25823 29121 25835 29155
rect 25777 29115 25835 29121
rect 25869 29155 25927 29161
rect 25869 29121 25881 29155
rect 25915 29121 25927 29155
rect 25869 29115 25927 29121
rect 25792 29084 25820 29115
rect 25958 29112 25964 29164
rect 26016 29152 26022 29164
rect 26344 29161 26372 29192
rect 26436 29192 26556 29220
rect 27264 29192 27384 29220
rect 27525 29223 27583 29229
rect 26436 29161 26464 29192
rect 26145 29155 26203 29161
rect 26145 29152 26157 29155
rect 26016 29124 26157 29152
rect 26016 29112 26022 29124
rect 26145 29121 26157 29124
rect 26191 29121 26203 29155
rect 26145 29115 26203 29121
rect 26329 29155 26387 29161
rect 26329 29121 26341 29155
rect 26375 29121 26387 29155
rect 26329 29115 26387 29121
rect 26421 29155 26479 29161
rect 26421 29121 26433 29155
rect 26467 29121 26479 29155
rect 26421 29115 26479 29121
rect 26513 29155 26571 29161
rect 26513 29121 26525 29155
rect 26559 29152 26571 29155
rect 26878 29152 26884 29164
rect 26559 29124 26884 29152
rect 26559 29121 26571 29124
rect 26513 29115 26571 29121
rect 26878 29112 26884 29124
rect 26936 29112 26942 29164
rect 27264 29161 27292 29192
rect 27525 29189 27537 29223
rect 27571 29220 27583 29223
rect 27908 29220 27936 29260
rect 28350 29248 28356 29260
rect 28408 29248 28414 29300
rect 28994 29248 29000 29300
rect 29052 29248 29058 29300
rect 29270 29248 29276 29300
rect 29328 29248 29334 29300
rect 30926 29248 30932 29300
rect 30984 29248 30990 29300
rect 31570 29248 31576 29300
rect 31628 29248 31634 29300
rect 31662 29248 31668 29300
rect 31720 29288 31726 29300
rect 31720 29260 32536 29288
rect 31720 29248 31726 29260
rect 29288 29220 29316 29248
rect 30834 29220 30840 29232
rect 27571 29192 27936 29220
rect 29196 29192 29316 29220
rect 30682 29192 30840 29220
rect 27571 29189 27583 29192
rect 27525 29183 27583 29189
rect 27249 29155 27307 29161
rect 27249 29121 27261 29155
rect 27295 29121 27307 29155
rect 27249 29115 27307 29121
rect 28626 29112 28632 29164
rect 28684 29112 28690 29164
rect 29196 29161 29224 29192
rect 30834 29180 30840 29192
rect 30892 29180 30898 29232
rect 30944 29220 30972 29248
rect 30944 29192 31800 29220
rect 29181 29155 29239 29161
rect 29181 29121 29193 29155
rect 29227 29121 29239 29155
rect 29181 29115 29239 29121
rect 31478 29112 31484 29164
rect 31536 29112 31542 29164
rect 31772 29161 31800 29192
rect 32508 29183 32536 29260
rect 34790 29248 34796 29300
rect 34848 29288 34854 29300
rect 34977 29291 35035 29297
rect 34977 29288 34989 29291
rect 34848 29260 34989 29288
rect 34848 29248 34854 29260
rect 34977 29257 34989 29260
rect 35023 29257 35035 29291
rect 34977 29251 35035 29257
rect 32494 29177 32552 29183
rect 34330 29180 34336 29232
rect 34388 29220 34394 29232
rect 34388 29192 35112 29220
rect 34388 29180 34394 29192
rect 31757 29155 31815 29161
rect 31757 29121 31769 29155
rect 31803 29121 31815 29155
rect 31757 29115 31815 29121
rect 31941 29155 31999 29161
rect 31941 29121 31953 29155
rect 31987 29152 31999 29155
rect 32125 29155 32183 29161
rect 32125 29152 32137 29155
rect 31987 29124 32137 29152
rect 31987 29121 31999 29124
rect 31941 29115 31999 29121
rect 32125 29121 32137 29124
rect 32171 29121 32183 29155
rect 32125 29115 32183 29121
rect 32306 29112 32312 29164
rect 32364 29112 32370 29164
rect 32401 29155 32459 29161
rect 32401 29121 32413 29155
rect 32447 29121 32459 29155
rect 32494 29143 32506 29177
rect 32540 29143 32552 29177
rect 32494 29137 32552 29143
rect 32401 29115 32459 29121
rect 30006 29084 30012 29096
rect 25792 29056 30012 29084
rect 30006 29044 30012 29056
rect 30064 29084 30070 29096
rect 30929 29087 30987 29093
rect 30929 29084 30941 29087
rect 30064 29056 30941 29084
rect 30064 29044 30070 29056
rect 30929 29053 30941 29056
rect 30975 29053 30987 29087
rect 32324 29084 32352 29112
rect 30929 29047 30987 29053
rect 31036 29056 32352 29084
rect 32416 29084 32444 29115
rect 33042 29112 33048 29164
rect 33100 29112 33106 29164
rect 34514 29112 34520 29164
rect 34572 29152 34578 29164
rect 34609 29155 34667 29161
rect 34609 29152 34621 29155
rect 34572 29124 34621 29152
rect 34572 29112 34578 29124
rect 34609 29121 34621 29124
rect 34655 29121 34667 29155
rect 34609 29115 34667 29121
rect 34974 29112 34980 29164
rect 35032 29112 35038 29164
rect 35084 29161 35112 29192
rect 35069 29155 35127 29161
rect 35069 29121 35081 29155
rect 35115 29121 35127 29155
rect 35069 29115 35127 29121
rect 36630 29112 36636 29164
rect 36688 29112 36694 29164
rect 36814 29112 36820 29164
rect 36872 29112 36878 29164
rect 33226 29084 33232 29096
rect 32416 29056 33232 29084
rect 26694 29016 26700 29028
rect 25516 28988 26700 29016
rect 26694 28976 26700 28988
rect 26752 28976 26758 29028
rect 26789 29019 26847 29025
rect 26789 28985 26801 29019
rect 26835 29016 26847 29019
rect 27062 29016 27068 29028
rect 26835 28988 27068 29016
rect 26835 28985 26847 28988
rect 26789 28979 26847 28985
rect 27062 28976 27068 28988
rect 27120 28976 27126 29028
rect 31036 29016 31064 29056
rect 30484 28988 31064 29016
rect 23400 28920 23612 28948
rect 24026 28908 24032 28960
rect 24084 28908 24090 28960
rect 25406 28908 25412 28960
rect 25464 28948 25470 28960
rect 25958 28948 25964 28960
rect 25464 28920 25964 28948
rect 25464 28908 25470 28920
rect 25958 28908 25964 28920
rect 26016 28908 26022 28960
rect 29270 28908 29276 28960
rect 29328 28948 29334 28960
rect 29438 28951 29496 28957
rect 29438 28948 29450 28951
rect 29328 28920 29450 28948
rect 29328 28908 29334 28920
rect 29438 28917 29450 28920
rect 29484 28917 29496 28951
rect 29438 28911 29496 28917
rect 30190 28908 30196 28960
rect 30248 28948 30254 28960
rect 30484 28948 30512 28988
rect 31110 28976 31116 29028
rect 31168 29016 31174 29028
rect 32416 29016 32444 29056
rect 33226 29044 33232 29056
rect 33284 29044 33290 29096
rect 31168 28988 32444 29016
rect 32769 29019 32827 29025
rect 31168 28976 31174 28988
rect 32769 28985 32781 29019
rect 32815 29016 32827 29019
rect 34698 29016 34704 29028
rect 32815 28988 34704 29016
rect 32815 28985 32827 28988
rect 32769 28979 32827 28985
rect 34698 28976 34704 28988
rect 34756 28976 34762 29028
rect 34793 29019 34851 29025
rect 34793 28985 34805 29019
rect 34839 29016 34851 29019
rect 34992 29016 35020 29112
rect 34839 28988 35020 29016
rect 37001 29019 37059 29025
rect 34839 28985 34851 28988
rect 34793 28979 34851 28985
rect 37001 28985 37013 29019
rect 37047 29016 37059 29019
rect 37274 29016 37280 29028
rect 37047 28988 37280 29016
rect 37047 28985 37059 28988
rect 37001 28979 37059 28985
rect 37274 28976 37280 28988
rect 37332 28976 37338 29028
rect 30248 28920 30512 28948
rect 30248 28908 30254 28920
rect 32398 28908 32404 28960
rect 32456 28948 32462 28960
rect 32861 28951 32919 28957
rect 32861 28948 32873 28951
rect 32456 28920 32873 28948
rect 32456 28908 32462 28920
rect 32861 28917 32873 28920
rect 32907 28917 32919 28951
rect 32861 28911 32919 28917
rect 1104 28858 38272 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38272 28858
rect 1104 28784 38272 28806
rect 4525 28747 4583 28753
rect 4525 28713 4537 28747
rect 4571 28744 4583 28747
rect 4614 28744 4620 28756
rect 4571 28716 4620 28744
rect 4571 28713 4583 28716
rect 4525 28707 4583 28713
rect 4614 28704 4620 28716
rect 4672 28704 4678 28756
rect 7929 28747 7987 28753
rect 7929 28713 7941 28747
rect 7975 28744 7987 28747
rect 8478 28744 8484 28756
rect 7975 28716 8484 28744
rect 7975 28713 7987 28716
rect 7929 28707 7987 28713
rect 8478 28704 8484 28716
rect 8536 28704 8542 28756
rect 20254 28744 20260 28756
rect 12406 28716 20260 28744
rect 5997 28611 6055 28617
rect 5997 28577 6009 28611
rect 6043 28608 6055 28611
rect 6181 28611 6239 28617
rect 6181 28608 6193 28611
rect 6043 28580 6193 28608
rect 6043 28577 6055 28580
rect 5997 28571 6055 28577
rect 6181 28577 6193 28580
rect 6227 28577 6239 28611
rect 6181 28571 6239 28577
rect 6457 28611 6515 28617
rect 6457 28577 6469 28611
rect 6503 28608 6515 28611
rect 6546 28608 6552 28620
rect 6503 28580 6552 28608
rect 6503 28577 6515 28580
rect 6457 28571 6515 28577
rect 6546 28568 6552 28580
rect 6604 28568 6610 28620
rect 12406 28608 12434 28716
rect 20254 28704 20260 28716
rect 20312 28704 20318 28756
rect 25590 28704 25596 28756
rect 25648 28744 25654 28756
rect 25777 28747 25835 28753
rect 25777 28744 25789 28747
rect 25648 28716 25789 28744
rect 25648 28704 25654 28716
rect 25777 28713 25789 28716
rect 25823 28713 25835 28747
rect 29086 28744 29092 28756
rect 25777 28707 25835 28713
rect 26252 28716 29092 28744
rect 16298 28636 16304 28688
rect 16356 28676 16362 28688
rect 26252 28676 26280 28716
rect 29086 28704 29092 28716
rect 29144 28704 29150 28756
rect 29270 28704 29276 28756
rect 29328 28704 29334 28756
rect 31588 28716 34008 28744
rect 31588 28688 31616 28716
rect 16356 28648 19334 28676
rect 16356 28636 16362 28648
rect 8312 28580 12434 28608
rect 16132 28580 18000 28608
rect 4341 28543 4399 28549
rect 4341 28509 4353 28543
rect 4387 28509 4399 28543
rect 4341 28503 4399 28509
rect 4709 28543 4767 28549
rect 4709 28509 4721 28543
rect 4755 28540 4767 28543
rect 5442 28540 5448 28552
rect 4755 28512 5448 28540
rect 4755 28509 4767 28512
rect 4709 28503 4767 28509
rect 4356 28472 4384 28503
rect 5442 28500 5448 28512
rect 5500 28500 5506 28552
rect 5626 28500 5632 28552
rect 5684 28500 5690 28552
rect 8312 28549 8340 28580
rect 16132 28552 16160 28580
rect 17972 28552 18000 28580
rect 18322 28568 18328 28620
rect 18380 28608 18386 28620
rect 18966 28608 18972 28620
rect 18380 28580 18972 28608
rect 18380 28568 18386 28580
rect 18966 28568 18972 28580
rect 19024 28568 19030 28620
rect 19306 28608 19334 28648
rect 19720 28648 21036 28676
rect 19610 28608 19616 28620
rect 19306 28580 19616 28608
rect 19610 28568 19616 28580
rect 19668 28568 19674 28620
rect 6089 28543 6147 28549
rect 6089 28509 6101 28543
rect 6135 28509 6147 28543
rect 6089 28503 6147 28509
rect 8297 28543 8355 28549
rect 8297 28509 8309 28543
rect 8343 28509 8355 28543
rect 8297 28503 8355 28509
rect 5644 28472 5672 28500
rect 4356 28444 5672 28472
rect 4246 28364 4252 28416
rect 4304 28364 4310 28416
rect 6104 28404 6132 28503
rect 7190 28432 7196 28484
rect 7248 28432 7254 28484
rect 8110 28472 8116 28484
rect 7760 28444 8116 28472
rect 7760 28404 7788 28444
rect 8110 28432 8116 28444
rect 8168 28472 8174 28484
rect 8312 28472 8340 28503
rect 9950 28500 9956 28552
rect 10008 28500 10014 28552
rect 10045 28543 10103 28549
rect 10045 28509 10057 28543
rect 10091 28540 10103 28543
rect 10229 28543 10287 28549
rect 10229 28540 10241 28543
rect 10091 28512 10241 28540
rect 10091 28509 10103 28512
rect 10045 28503 10103 28509
rect 10229 28509 10241 28512
rect 10275 28509 10287 28543
rect 10229 28503 10287 28509
rect 13446 28500 13452 28552
rect 13504 28540 13510 28552
rect 14274 28540 14280 28552
rect 13504 28512 14280 28540
rect 13504 28500 13510 28512
rect 14274 28500 14280 28512
rect 14332 28500 14338 28552
rect 16114 28500 16120 28552
rect 16172 28500 16178 28552
rect 16206 28500 16212 28552
rect 16264 28540 16270 28552
rect 16301 28543 16359 28549
rect 16301 28540 16313 28543
rect 16264 28512 16313 28540
rect 16264 28500 16270 28512
rect 16301 28509 16313 28512
rect 16347 28509 16359 28543
rect 16301 28503 16359 28509
rect 16482 28500 16488 28552
rect 16540 28500 16546 28552
rect 17954 28500 17960 28552
rect 18012 28500 18018 28552
rect 19720 28549 19748 28648
rect 19886 28568 19892 28620
rect 19944 28608 19950 28620
rect 19944 28580 20116 28608
rect 19944 28568 19950 28580
rect 20088 28549 20116 28580
rect 21008 28552 21036 28648
rect 24872 28648 26280 28676
rect 24486 28608 24492 28620
rect 22388 28580 24492 28608
rect 22388 28552 22416 28580
rect 24486 28568 24492 28580
rect 24544 28608 24550 28620
rect 24544 28580 24624 28608
rect 24544 28568 24550 28580
rect 19705 28543 19763 28549
rect 19705 28540 19717 28543
rect 19276 28512 19717 28540
rect 8168 28444 8340 28472
rect 9968 28472 9996 28500
rect 10410 28472 10416 28484
rect 9968 28444 10416 28472
rect 8168 28432 8174 28444
rect 10410 28432 10416 28444
rect 10468 28432 10474 28484
rect 10502 28432 10508 28484
rect 10560 28432 10566 28484
rect 11054 28432 11060 28484
rect 11112 28432 11118 28484
rect 14090 28472 14096 28484
rect 11992 28444 14096 28472
rect 11992 28416 12020 28444
rect 14090 28432 14096 28444
rect 14148 28472 14154 28484
rect 16393 28475 16451 28481
rect 16393 28472 16405 28475
rect 14148 28444 16405 28472
rect 14148 28432 14154 28444
rect 16393 28441 16405 28444
rect 16439 28472 16451 28475
rect 16850 28472 16856 28484
rect 16439 28444 16856 28472
rect 16439 28441 16451 28444
rect 16393 28435 16451 28441
rect 16850 28432 16856 28444
rect 16908 28432 16914 28484
rect 17862 28432 17868 28484
rect 17920 28472 17926 28484
rect 19276 28472 19304 28512
rect 19705 28509 19717 28512
rect 19751 28509 19763 28543
rect 19705 28503 19763 28509
rect 19797 28543 19855 28549
rect 19797 28509 19809 28543
rect 19843 28540 19855 28543
rect 20073 28543 20131 28549
rect 19843 28512 20024 28540
rect 19843 28509 19855 28512
rect 19797 28503 19855 28509
rect 17920 28444 19304 28472
rect 17920 28432 17926 28444
rect 19334 28432 19340 28484
rect 19392 28472 19398 28484
rect 19889 28475 19947 28481
rect 19889 28472 19901 28475
rect 19392 28444 19901 28472
rect 19392 28432 19398 28444
rect 19889 28441 19901 28444
rect 19935 28441 19947 28475
rect 19996 28472 20024 28512
rect 20073 28509 20085 28543
rect 20119 28509 20131 28543
rect 20073 28503 20131 28509
rect 20622 28500 20628 28552
rect 20680 28500 20686 28552
rect 20806 28500 20812 28552
rect 20864 28500 20870 28552
rect 20990 28500 20996 28552
rect 21048 28500 21054 28552
rect 21266 28500 21272 28552
rect 21324 28540 21330 28552
rect 21634 28540 21640 28552
rect 21324 28512 21640 28540
rect 21324 28500 21330 28512
rect 21634 28500 21640 28512
rect 21692 28500 21698 28552
rect 22002 28500 22008 28552
rect 22060 28500 22066 28552
rect 22370 28500 22376 28552
rect 22428 28500 22434 28552
rect 22465 28543 22523 28549
rect 22465 28509 22477 28543
rect 22511 28540 22523 28543
rect 22554 28540 22560 28552
rect 22511 28512 22560 28540
rect 22511 28509 22523 28512
rect 22465 28503 22523 28509
rect 22554 28500 22560 28512
rect 22612 28500 22618 28552
rect 22922 28500 22928 28552
rect 22980 28540 22986 28552
rect 23750 28540 23756 28552
rect 22980 28512 23756 28540
rect 22980 28500 22986 28512
rect 23750 28500 23756 28512
rect 23808 28500 23814 28552
rect 24596 28549 24624 28580
rect 24581 28543 24639 28549
rect 24581 28509 24593 28543
rect 24627 28509 24639 28543
rect 24581 28503 24639 28509
rect 24670 28500 24676 28552
rect 24728 28540 24734 28552
rect 24872 28540 24900 28648
rect 26142 28608 26148 28620
rect 25976 28580 26148 28608
rect 24728 28512 24900 28540
rect 24728 28500 24734 28512
rect 24946 28500 24952 28552
rect 25004 28500 25010 28552
rect 25314 28500 25320 28552
rect 25372 28500 25378 28552
rect 25590 28500 25596 28552
rect 25648 28540 25654 28552
rect 25976 28549 26004 28580
rect 26142 28568 26148 28580
rect 26200 28568 26206 28620
rect 25961 28543 26019 28549
rect 25961 28540 25973 28543
rect 25648 28512 25973 28540
rect 25648 28500 25654 28512
rect 25961 28509 25973 28512
rect 26007 28509 26019 28543
rect 25961 28503 26019 28509
rect 26053 28543 26111 28549
rect 26053 28509 26065 28543
rect 26099 28540 26111 28543
rect 26252 28540 26280 28648
rect 26344 28648 30788 28676
rect 26344 28549 26372 28648
rect 30006 28568 30012 28620
rect 30064 28568 30070 28620
rect 30098 28568 30104 28620
rect 30156 28568 30162 28620
rect 30760 28608 30788 28648
rect 31570 28636 31576 28688
rect 31628 28636 31634 28688
rect 33980 28676 34008 28716
rect 33980 28648 34100 28676
rect 32033 28611 32091 28617
rect 30760 28580 31708 28608
rect 26099 28512 26280 28540
rect 26329 28543 26387 28549
rect 26099 28509 26111 28512
rect 26053 28503 26111 28509
rect 26329 28509 26341 28543
rect 26375 28509 26387 28543
rect 26329 28503 26387 28509
rect 29089 28543 29147 28549
rect 29089 28509 29101 28543
rect 29135 28540 29147 28543
rect 29135 28512 29592 28540
rect 29135 28509 29147 28512
rect 29089 28503 29147 28509
rect 20640 28472 20668 28500
rect 19996 28444 20668 28472
rect 22020 28472 22048 28500
rect 22020 28444 24716 28472
rect 19889 28435 19947 28441
rect 6104 28376 7788 28404
rect 7926 28364 7932 28416
rect 7984 28404 7990 28416
rect 8205 28407 8263 28413
rect 8205 28404 8217 28407
rect 7984 28376 8217 28404
rect 7984 28364 7990 28376
rect 8205 28373 8217 28376
rect 8251 28373 8263 28407
rect 8205 28367 8263 28373
rect 11974 28364 11980 28416
rect 12032 28364 12038 28416
rect 16482 28364 16488 28416
rect 16540 28404 16546 28416
rect 16669 28407 16727 28413
rect 16669 28404 16681 28407
rect 16540 28376 16681 28404
rect 16540 28364 16546 28376
rect 16669 28373 16681 28376
rect 16715 28373 16727 28407
rect 16669 28367 16727 28373
rect 19426 28364 19432 28416
rect 19484 28404 19490 28416
rect 19521 28407 19579 28413
rect 19521 28404 19533 28407
rect 19484 28376 19533 28404
rect 19484 28364 19490 28376
rect 19521 28373 19533 28376
rect 19567 28373 19579 28407
rect 19521 28367 19579 28373
rect 20162 28364 20168 28416
rect 20220 28404 20226 28416
rect 21082 28404 21088 28416
rect 20220 28376 21088 28404
rect 20220 28364 20226 28376
rect 21082 28364 21088 28376
rect 21140 28364 21146 28416
rect 21542 28364 21548 28416
rect 21600 28404 21606 28416
rect 23750 28404 23756 28416
rect 21600 28376 23756 28404
rect 21600 28364 21606 28376
rect 23750 28364 23756 28376
rect 23808 28364 23814 28416
rect 24394 28364 24400 28416
rect 24452 28364 24458 28416
rect 24688 28404 24716 28444
rect 24762 28432 24768 28484
rect 24820 28432 24826 28484
rect 25332 28472 25360 28500
rect 25866 28472 25872 28484
rect 25332 28444 25872 28472
rect 25866 28432 25872 28444
rect 25924 28472 25930 28484
rect 26145 28475 26203 28481
rect 26145 28472 26157 28475
rect 25924 28444 26157 28472
rect 25924 28432 25930 28444
rect 26145 28441 26157 28444
rect 26191 28441 26203 28475
rect 26145 28435 26203 28441
rect 24946 28404 24952 28416
rect 24688 28376 24952 28404
rect 24946 28364 24952 28376
rect 25004 28404 25010 28416
rect 26344 28404 26372 28503
rect 29564 28413 29592 28512
rect 30024 28472 30052 28568
rect 30374 28500 30380 28552
rect 30432 28500 30438 28552
rect 30760 28549 30788 28580
rect 30470 28543 30528 28549
rect 30470 28509 30482 28543
rect 30516 28509 30528 28543
rect 30470 28503 30528 28509
rect 30745 28543 30803 28549
rect 30745 28509 30757 28543
rect 30791 28509 30803 28543
rect 30745 28503 30803 28509
rect 30842 28543 30900 28549
rect 30842 28509 30854 28543
rect 30888 28540 30900 28543
rect 31297 28543 31355 28549
rect 31297 28540 31309 28543
rect 30888 28512 30972 28540
rect 30888 28509 30900 28512
rect 30842 28503 30900 28509
rect 30484 28472 30512 28503
rect 30024 28444 30512 28472
rect 30650 28432 30656 28484
rect 30708 28432 30714 28484
rect 30944 28416 30972 28512
rect 31036 28512 31309 28540
rect 25004 28376 26372 28404
rect 29549 28407 29607 28413
rect 25004 28364 25010 28376
rect 29549 28373 29561 28407
rect 29595 28373 29607 28407
rect 29549 28367 29607 28373
rect 29917 28407 29975 28413
rect 29917 28373 29929 28407
rect 29963 28404 29975 28407
rect 30190 28404 30196 28416
rect 29963 28376 30196 28404
rect 29963 28373 29975 28376
rect 29917 28367 29975 28373
rect 30190 28364 30196 28376
rect 30248 28364 30254 28416
rect 30926 28364 30932 28416
rect 30984 28364 30990 28416
rect 31036 28413 31064 28512
rect 31297 28509 31309 28512
rect 31343 28509 31355 28543
rect 31297 28503 31355 28509
rect 31478 28500 31484 28552
rect 31536 28540 31542 28552
rect 31573 28543 31631 28549
rect 31573 28540 31585 28543
rect 31536 28512 31585 28540
rect 31536 28500 31542 28512
rect 31573 28509 31585 28512
rect 31619 28509 31631 28543
rect 31573 28503 31631 28509
rect 31680 28472 31708 28580
rect 32033 28577 32045 28611
rect 32079 28608 32091 28611
rect 32398 28608 32404 28620
rect 32079 28580 32404 28608
rect 32079 28577 32091 28580
rect 32033 28571 32091 28577
rect 32398 28568 32404 28580
rect 32456 28568 32462 28620
rect 33318 28568 33324 28620
rect 33376 28608 33382 28620
rect 33873 28611 33931 28617
rect 33873 28608 33885 28611
rect 33376 28580 33885 28608
rect 33376 28568 33382 28580
rect 33873 28577 33885 28580
rect 33919 28608 33931 28611
rect 33962 28608 33968 28620
rect 33919 28580 33968 28608
rect 33919 28577 33931 28580
rect 33873 28571 33931 28577
rect 33962 28568 33968 28580
rect 34020 28568 34026 28620
rect 34072 28617 34100 28648
rect 34057 28611 34115 28617
rect 34057 28577 34069 28611
rect 34103 28608 34115 28611
rect 36449 28611 36507 28617
rect 36449 28608 36461 28611
rect 34103 28580 36461 28608
rect 34103 28577 34115 28580
rect 34057 28571 34115 28577
rect 36449 28577 36461 28580
rect 36495 28577 36507 28611
rect 36449 28571 36507 28577
rect 31754 28500 31760 28552
rect 31812 28500 31818 28552
rect 34698 28500 34704 28552
rect 34756 28500 34762 28552
rect 31938 28472 31944 28484
rect 31680 28444 31944 28472
rect 31938 28432 31944 28444
rect 31996 28432 32002 28484
rect 34054 28472 34060 28484
rect 33258 28444 34060 28472
rect 34054 28432 34060 28444
rect 34112 28432 34118 28484
rect 34422 28432 34428 28484
rect 34480 28472 34486 28484
rect 34977 28475 35035 28481
rect 34977 28472 34989 28475
rect 34480 28444 34989 28472
rect 34480 28432 34486 28444
rect 34977 28441 34989 28444
rect 35023 28441 35035 28475
rect 34977 28435 35035 28441
rect 35986 28432 35992 28484
rect 36044 28432 36050 28484
rect 31021 28407 31079 28413
rect 31021 28373 31033 28407
rect 31067 28373 31079 28407
rect 31021 28367 31079 28373
rect 31110 28364 31116 28416
rect 31168 28364 31174 28416
rect 31478 28364 31484 28416
rect 31536 28364 31542 28416
rect 31956 28404 31984 28432
rect 33505 28407 33563 28413
rect 33505 28404 33517 28407
rect 31956 28376 33517 28404
rect 33505 28373 33517 28376
rect 33551 28373 33563 28407
rect 33505 28367 33563 28373
rect 34146 28364 34152 28416
rect 34204 28364 34210 28416
rect 34514 28364 34520 28416
rect 34572 28364 34578 28416
rect 1104 28314 38272 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38272 28314
rect 1104 28240 38272 28262
rect 4246 28160 4252 28212
rect 4304 28160 4310 28212
rect 6822 28160 6828 28212
rect 6880 28160 6886 28212
rect 9674 28200 9680 28212
rect 7208 28172 8248 28200
rect 4264 28132 4292 28160
rect 7208 28144 7236 28172
rect 4080 28104 4292 28132
rect 4341 28135 4399 28141
rect 4080 28073 4108 28104
rect 4341 28101 4353 28135
rect 4387 28132 4399 28135
rect 4614 28132 4620 28144
rect 4387 28104 4620 28132
rect 4387 28101 4399 28104
rect 4341 28095 4399 28101
rect 4614 28092 4620 28104
rect 4672 28092 4678 28144
rect 7190 28092 7196 28144
rect 7248 28092 7254 28144
rect 7926 28132 7932 28144
rect 7668 28104 7932 28132
rect 4065 28067 4123 28073
rect 4065 28033 4077 28067
rect 4111 28033 4123 28067
rect 4065 28027 4123 28033
rect 5350 28024 5356 28076
rect 5408 28064 5414 28076
rect 5994 28064 6000 28076
rect 5408 28036 6000 28064
rect 5408 28024 5414 28036
rect 5994 28024 6000 28036
rect 6052 28024 6058 28076
rect 7668 28073 7696 28104
rect 7926 28092 7932 28104
rect 7984 28092 7990 28144
rect 8220 28132 8248 28172
rect 8312 28172 9680 28200
rect 8312 28132 8340 28172
rect 9674 28160 9680 28172
rect 9732 28160 9738 28212
rect 10502 28160 10508 28212
rect 10560 28200 10566 28212
rect 10597 28203 10655 28209
rect 10597 28200 10609 28203
rect 10560 28172 10609 28200
rect 10560 28160 10566 28172
rect 10597 28169 10609 28172
rect 10643 28169 10655 28203
rect 10597 28163 10655 28169
rect 11517 28203 11575 28209
rect 11517 28169 11529 28203
rect 11563 28169 11575 28203
rect 11517 28163 11575 28169
rect 11885 28203 11943 28209
rect 11885 28169 11897 28203
rect 11931 28200 11943 28203
rect 11974 28200 11980 28212
rect 11931 28172 11980 28200
rect 11931 28169 11943 28172
rect 11885 28163 11943 28169
rect 8220 28104 8418 28132
rect 6733 28067 6791 28073
rect 6733 28033 6745 28067
rect 6779 28064 6791 28067
rect 7653 28067 7711 28073
rect 6779 28036 7604 28064
rect 6779 28033 6791 28036
rect 6733 28027 6791 28033
rect 5813 27999 5871 28005
rect 5813 27965 5825 27999
rect 5859 27996 5871 27999
rect 6748 27996 6776 28027
rect 5859 27968 6776 27996
rect 7009 27999 7067 28005
rect 5859 27965 5871 27968
rect 5813 27959 5871 27965
rect 7009 27965 7021 27999
rect 7055 27996 7067 27999
rect 7466 27996 7472 28008
rect 7055 27968 7472 27996
rect 7055 27965 7067 27968
rect 7009 27959 7067 27965
rect 7466 27956 7472 27968
rect 7524 27956 7530 28008
rect 6362 27820 6368 27872
rect 6420 27820 6426 27872
rect 7576 27860 7604 28036
rect 7653 28033 7665 28067
rect 7699 28033 7711 28067
rect 7653 28027 7711 28033
rect 9766 28024 9772 28076
rect 9824 28064 9830 28076
rect 9953 28067 10011 28073
rect 9953 28064 9965 28067
rect 9824 28036 9965 28064
rect 9824 28024 9830 28036
rect 9953 28033 9965 28036
rect 9999 28064 10011 28067
rect 10781 28067 10839 28073
rect 9999 28036 10732 28064
rect 9999 28033 10011 28036
rect 9953 28027 10011 28033
rect 7929 27999 7987 28005
rect 7929 27965 7941 27999
rect 7975 27996 7987 27999
rect 8294 27996 8300 28008
rect 7975 27968 8300 27996
rect 7975 27965 7987 27968
rect 7929 27959 7987 27965
rect 8294 27956 8300 27968
rect 8352 27956 8358 28008
rect 9401 27999 9459 28005
rect 9401 27965 9413 27999
rect 9447 27996 9459 27999
rect 10045 27999 10103 28005
rect 10045 27996 10057 27999
rect 9447 27968 10057 27996
rect 9447 27965 9459 27968
rect 9401 27959 9459 27965
rect 10045 27965 10057 27968
rect 10091 27965 10103 27999
rect 10045 27959 10103 27965
rect 10060 27928 10088 27959
rect 10134 27956 10140 28008
rect 10192 27956 10198 28008
rect 10704 27996 10732 28036
rect 10781 28033 10793 28067
rect 10827 28064 10839 28067
rect 11532 28064 11560 28163
rect 11974 28160 11980 28172
rect 12032 28200 12038 28212
rect 12032 28172 12480 28200
rect 12032 28160 12038 28172
rect 10827 28036 11560 28064
rect 12452 28073 12480 28172
rect 12526 28160 12532 28212
rect 12584 28160 12590 28212
rect 13446 28160 13452 28212
rect 13504 28200 13510 28212
rect 13725 28203 13783 28209
rect 13725 28200 13737 28203
rect 13504 28172 13737 28200
rect 13504 28160 13510 28172
rect 13725 28169 13737 28172
rect 13771 28169 13783 28203
rect 13725 28163 13783 28169
rect 13909 28203 13967 28209
rect 13909 28169 13921 28203
rect 13955 28200 13967 28203
rect 13998 28200 14004 28212
rect 13955 28172 14004 28200
rect 13955 28169 13967 28172
rect 13909 28163 13967 28169
rect 13998 28160 14004 28172
rect 14056 28160 14062 28212
rect 14829 28203 14887 28209
rect 14829 28169 14841 28203
rect 14875 28200 14887 28203
rect 16114 28200 16120 28212
rect 14875 28172 16120 28200
rect 14875 28169 14887 28172
rect 14829 28163 14887 28169
rect 16114 28160 16120 28172
rect 16172 28160 16178 28212
rect 16574 28160 16580 28212
rect 16632 28200 16638 28212
rect 16632 28172 18000 28200
rect 16632 28160 16638 28172
rect 12544 28132 12572 28160
rect 12621 28135 12679 28141
rect 12621 28132 12633 28135
rect 12544 28104 12633 28132
rect 12621 28101 12633 28104
rect 12667 28101 12679 28135
rect 14016 28132 14044 28160
rect 15838 28132 15844 28144
rect 14016 28104 15844 28132
rect 12621 28095 12679 28101
rect 15838 28092 15844 28104
rect 15896 28092 15902 28144
rect 16850 28092 16856 28144
rect 16908 28132 16914 28144
rect 17037 28135 17095 28141
rect 17037 28132 17049 28135
rect 16908 28104 17049 28132
rect 16908 28092 16914 28104
rect 17037 28101 17049 28104
rect 17083 28101 17095 28135
rect 17037 28095 17095 28101
rect 12452 28067 12515 28073
rect 12452 28036 12469 28067
rect 10827 28033 10839 28036
rect 10781 28027 10839 28033
rect 12457 28033 12469 28036
rect 12503 28033 12515 28067
rect 12457 28027 12515 28033
rect 12713 28067 12771 28073
rect 12713 28033 12725 28067
rect 12759 28033 12771 28067
rect 12713 28027 12771 28033
rect 12805 28067 12863 28073
rect 12805 28033 12817 28067
rect 12851 28064 12863 28067
rect 13170 28064 13176 28076
rect 12851 28036 13176 28064
rect 12851 28033 12863 28036
rect 12805 28027 12863 28033
rect 11974 27996 11980 28008
rect 10704 27968 11980 27996
rect 11974 27956 11980 27968
rect 12032 27956 12038 28008
rect 12066 27956 12072 28008
rect 12124 27956 12130 28008
rect 12728 27996 12756 28027
rect 13170 28024 13176 28036
rect 13228 28024 13234 28076
rect 13817 28067 13875 28073
rect 13817 28033 13829 28067
rect 13863 28064 13875 28067
rect 14366 28064 14372 28076
rect 13863 28036 14372 28064
rect 13863 28033 13875 28036
rect 13817 28027 13875 28033
rect 14366 28024 14372 28036
rect 14424 28024 14430 28076
rect 14550 28024 14556 28076
rect 14608 28064 14614 28076
rect 14921 28067 14979 28073
rect 14921 28064 14933 28067
rect 14608 28036 14933 28064
rect 14608 28024 14614 28036
rect 14921 28033 14933 28036
rect 14967 28064 14979 28067
rect 15194 28064 15200 28076
rect 14967 28036 15200 28064
rect 14967 28033 14979 28036
rect 14921 28027 14979 28033
rect 15194 28024 15200 28036
rect 15252 28024 15258 28076
rect 16022 28024 16028 28076
rect 16080 28064 16086 28076
rect 16669 28067 16727 28073
rect 16669 28064 16681 28067
rect 16080 28036 16681 28064
rect 16080 28024 16086 28036
rect 16669 28033 16681 28036
rect 16715 28033 16727 28067
rect 16669 28027 16727 28033
rect 16758 28024 16764 28076
rect 16816 28064 16822 28076
rect 16945 28067 17003 28073
rect 16816 28036 16861 28064
rect 16816 28024 16822 28036
rect 16945 28033 16957 28067
rect 16991 28033 17003 28067
rect 16945 28027 17003 28033
rect 17175 28067 17233 28073
rect 17175 28033 17187 28067
rect 17221 28064 17233 28067
rect 17310 28064 17316 28076
rect 17221 28036 17316 28064
rect 17221 28033 17233 28036
rect 17175 28027 17233 28033
rect 13541 27999 13599 28005
rect 13541 27996 13553 27999
rect 12728 27968 13553 27996
rect 12728 27928 12756 27968
rect 13541 27965 13553 27968
rect 13587 27996 13599 27999
rect 16776 27996 16804 28024
rect 13587 27968 16804 27996
rect 16960 27996 16988 28027
rect 17310 28024 17316 28036
rect 17368 28064 17374 28076
rect 17862 28064 17868 28076
rect 17368 28036 17868 28064
rect 17368 28024 17374 28036
rect 17862 28024 17868 28036
rect 17920 28024 17926 28076
rect 17972 28064 18000 28172
rect 18414 28160 18420 28212
rect 18472 28160 18478 28212
rect 18782 28160 18788 28212
rect 18840 28200 18846 28212
rect 18840 28172 19196 28200
rect 18840 28160 18846 28172
rect 18432 28132 18460 28160
rect 19168 28144 19196 28172
rect 19536 28172 21220 28200
rect 19061 28135 19119 28141
rect 19061 28132 19073 28135
rect 18432 28104 19073 28132
rect 19061 28101 19073 28104
rect 19107 28101 19119 28135
rect 19061 28095 19119 28101
rect 18782 28064 18788 28076
rect 17972 28036 18788 28064
rect 18782 28024 18788 28036
rect 18840 28024 18846 28076
rect 19076 28064 19104 28095
rect 19150 28092 19156 28144
rect 19208 28132 19214 28144
rect 19261 28135 19319 28141
rect 19261 28132 19273 28135
rect 19208 28104 19273 28132
rect 19208 28092 19214 28104
rect 19261 28101 19273 28104
rect 19307 28101 19319 28135
rect 19261 28095 19319 28101
rect 19536 28064 19564 28172
rect 20714 28132 20720 28144
rect 19628 28104 20720 28132
rect 19628 28073 19656 28104
rect 20714 28092 20720 28104
rect 20772 28092 20778 28144
rect 21192 28132 21220 28172
rect 21284 28172 21404 28200
rect 21284 28132 21312 28172
rect 20824 28104 21036 28132
rect 19076 28036 19564 28064
rect 19613 28067 19671 28073
rect 19613 28033 19625 28067
rect 19659 28033 19671 28067
rect 19899 28067 19957 28073
rect 19899 28042 19911 28067
rect 19613 28027 19671 28033
rect 19334 27996 19340 28008
rect 16960 27968 19340 27996
rect 13587 27965 13599 27968
rect 13541 27959 13599 27965
rect 19334 27956 19340 27968
rect 19392 27956 19398 28008
rect 19518 27956 19524 28008
rect 19576 27996 19582 28008
rect 19797 27999 19855 28005
rect 19797 27996 19809 27999
rect 19576 27968 19809 27996
rect 19576 27956 19582 27968
rect 19797 27965 19809 27968
rect 19843 27965 19855 27999
rect 19886 27990 19892 28042
rect 19945 28033 19957 28067
rect 19944 28027 19957 28033
rect 19944 27990 19950 28027
rect 20070 28024 20076 28076
rect 20128 28024 20134 28076
rect 20824 28073 20852 28104
rect 20625 28067 20683 28073
rect 20625 28033 20637 28067
rect 20671 28064 20683 28067
rect 20809 28067 20867 28073
rect 20809 28064 20821 28067
rect 20671 28036 20821 28064
rect 20671 28033 20683 28036
rect 20625 28027 20683 28033
rect 20809 28033 20821 28036
rect 20855 28033 20867 28067
rect 20809 28027 20867 28033
rect 20902 28067 20960 28073
rect 20902 28033 20914 28067
rect 20948 28033 20960 28067
rect 20902 28027 20960 28033
rect 20165 27999 20223 28005
rect 20165 27996 20177 27999
rect 19797 27959 19855 27965
rect 19996 27968 20177 27996
rect 8956 27900 9720 27928
rect 10060 27900 12756 27928
rect 14093 27931 14151 27937
rect 8956 27860 8984 27900
rect 9692 27872 9720 27900
rect 14093 27897 14105 27931
rect 14139 27928 14151 27931
rect 14553 27931 14611 27937
rect 14553 27928 14565 27931
rect 14139 27900 14565 27928
rect 14139 27897 14151 27900
rect 14093 27891 14151 27897
rect 14553 27897 14565 27900
rect 14599 27897 14611 27931
rect 14553 27891 14611 27897
rect 14642 27888 14648 27940
rect 14700 27888 14706 27940
rect 15746 27888 15752 27940
rect 15804 27928 15810 27940
rect 19429 27931 19487 27937
rect 15804 27900 19288 27928
rect 15804 27888 15810 27900
rect 16132 27872 16160 27900
rect 7576 27832 8984 27860
rect 9490 27820 9496 27872
rect 9548 27860 9554 27872
rect 9585 27863 9643 27869
rect 9585 27860 9597 27863
rect 9548 27832 9597 27860
rect 9548 27820 9554 27832
rect 9585 27829 9597 27832
rect 9631 27829 9643 27863
rect 9585 27823 9643 27829
rect 9674 27820 9680 27872
rect 9732 27820 9738 27872
rect 10962 27820 10968 27872
rect 11020 27860 11026 27872
rect 12066 27860 12072 27872
rect 11020 27832 12072 27860
rect 11020 27820 11026 27832
rect 12066 27820 12072 27832
rect 12124 27820 12130 27872
rect 12989 27863 13047 27869
rect 12989 27829 13001 27863
rect 13035 27860 13047 27863
rect 13630 27860 13636 27872
rect 13035 27832 13636 27860
rect 13035 27829 13047 27832
rect 12989 27823 13047 27829
rect 13630 27820 13636 27832
rect 13688 27820 13694 27872
rect 14182 27820 14188 27872
rect 14240 27820 14246 27872
rect 14458 27820 14464 27872
rect 14516 27860 14522 27872
rect 15470 27860 15476 27872
rect 14516 27832 15476 27860
rect 14516 27820 14522 27832
rect 15470 27820 15476 27832
rect 15528 27820 15534 27872
rect 16114 27820 16120 27872
rect 16172 27820 16178 27872
rect 17310 27820 17316 27872
rect 17368 27820 17374 27872
rect 17402 27820 17408 27872
rect 17460 27860 17466 27872
rect 17678 27860 17684 27872
rect 17460 27832 17684 27860
rect 17460 27820 17466 27832
rect 17678 27820 17684 27832
rect 17736 27860 17742 27872
rect 18230 27860 18236 27872
rect 17736 27832 18236 27860
rect 17736 27820 17742 27832
rect 18230 27820 18236 27832
rect 18288 27820 18294 27872
rect 19260 27869 19288 27900
rect 19429 27897 19441 27931
rect 19475 27928 19487 27931
rect 19610 27928 19616 27940
rect 19475 27900 19616 27928
rect 19475 27897 19487 27900
rect 19429 27891 19487 27897
rect 19610 27888 19616 27900
rect 19668 27888 19674 27940
rect 19705 27931 19763 27937
rect 19705 27897 19717 27931
rect 19751 27928 19763 27931
rect 19996 27928 20024 27968
rect 20165 27965 20177 27968
rect 20211 27965 20223 27999
rect 20165 27959 20223 27965
rect 20346 27956 20352 28008
rect 20404 27956 20410 28008
rect 20441 27999 20499 28005
rect 20441 27965 20453 27999
rect 20487 27965 20499 27999
rect 20441 27959 20499 27965
rect 20533 27999 20591 28005
rect 20533 27965 20545 27999
rect 20579 27996 20591 27999
rect 20917 27996 20945 28027
rect 20579 27968 20945 27996
rect 20579 27965 20591 27968
rect 20533 27959 20591 27965
rect 19751 27900 20024 27928
rect 19751 27897 19763 27900
rect 19705 27891 19763 27897
rect 19245 27863 19303 27869
rect 19245 27829 19257 27863
rect 19291 27860 19303 27863
rect 19886 27860 19892 27872
rect 19291 27832 19892 27860
rect 19291 27829 19303 27832
rect 19245 27823 19303 27829
rect 19886 27820 19892 27832
rect 19944 27860 19950 27872
rect 20456 27860 20484 27959
rect 19944 27832 20484 27860
rect 19944 27820 19950 27832
rect 20530 27820 20536 27872
rect 20588 27860 20594 27872
rect 20732 27860 20760 27968
rect 21008 27928 21036 28104
rect 21192 28104 21312 28132
rect 21376 28132 21404 28172
rect 23014 28160 23020 28212
rect 23072 28200 23078 28212
rect 23109 28203 23167 28209
rect 23109 28200 23121 28203
rect 23072 28172 23121 28200
rect 23072 28160 23078 28172
rect 23109 28169 23121 28172
rect 23155 28169 23167 28203
rect 23109 28163 23167 28169
rect 23290 28160 23296 28212
rect 23348 28200 23354 28212
rect 23845 28203 23903 28209
rect 23845 28200 23857 28203
rect 23348 28172 23857 28200
rect 23348 28160 23354 28172
rect 23845 28169 23857 28172
rect 23891 28169 23903 28203
rect 23845 28163 23903 28169
rect 24210 28160 24216 28212
rect 24268 28200 24274 28212
rect 26786 28200 26792 28212
rect 24268 28172 26792 28200
rect 24268 28160 24274 28172
rect 26786 28160 26792 28172
rect 26844 28160 26850 28212
rect 29086 28160 29092 28212
rect 29144 28200 29150 28212
rect 31478 28200 31484 28212
rect 29144 28172 31484 28200
rect 29144 28160 29150 28172
rect 31478 28160 31484 28172
rect 31536 28160 31542 28212
rect 31754 28160 31760 28212
rect 31812 28200 31818 28212
rect 31849 28203 31907 28209
rect 31849 28200 31861 28203
rect 31812 28172 31861 28200
rect 31812 28160 31818 28172
rect 31849 28169 31861 28172
rect 31895 28169 31907 28203
rect 31849 28163 31907 28169
rect 31938 28160 31944 28212
rect 31996 28200 32002 28212
rect 32585 28203 32643 28209
rect 32585 28200 32597 28203
rect 31996 28172 32597 28200
rect 31996 28160 32002 28172
rect 32585 28169 32597 28172
rect 32631 28169 32643 28203
rect 32585 28163 32643 28169
rect 32953 28203 33011 28209
rect 32953 28169 32965 28203
rect 32999 28200 33011 28203
rect 33042 28200 33048 28212
rect 32999 28172 33048 28200
rect 32999 28169 33011 28172
rect 32953 28163 33011 28169
rect 33042 28160 33048 28172
rect 33100 28160 33106 28212
rect 34422 28160 34428 28212
rect 34480 28160 34486 28212
rect 34606 28160 34612 28212
rect 34664 28160 34670 28212
rect 34698 28160 34704 28212
rect 34756 28200 34762 28212
rect 34885 28203 34943 28209
rect 34885 28200 34897 28203
rect 34756 28172 34897 28200
rect 34756 28160 34762 28172
rect 34885 28169 34897 28172
rect 34931 28169 34943 28203
rect 34885 28163 34943 28169
rect 37274 28160 37280 28212
rect 37332 28160 37338 28212
rect 22186 28132 22192 28144
rect 21376 28104 22192 28132
rect 21192 28073 21220 28104
rect 22186 28092 22192 28104
rect 22244 28092 22250 28144
rect 34624 28132 34652 28160
rect 23676 28104 24716 28132
rect 21085 28067 21143 28073
rect 21085 28033 21097 28067
rect 21131 28033 21143 28067
rect 21085 28027 21143 28033
rect 21177 28067 21235 28073
rect 21177 28033 21189 28067
rect 21223 28033 21235 28067
rect 21177 28027 21235 28033
rect 21274 28067 21332 28073
rect 21274 28033 21286 28067
rect 21320 28064 21332 28067
rect 21450 28064 21456 28076
rect 21320 28036 21456 28064
rect 21320 28033 21332 28036
rect 21274 28027 21332 28033
rect 21100 27996 21128 28027
rect 21450 28024 21456 28036
rect 21508 28024 21514 28076
rect 21634 28024 21640 28076
rect 21692 28064 21698 28076
rect 22465 28067 22523 28073
rect 22465 28064 22477 28067
rect 21692 28036 22477 28064
rect 21692 28024 21698 28036
rect 22465 28033 22477 28036
rect 22511 28033 22523 28067
rect 22465 28027 22523 28033
rect 22833 28067 22891 28073
rect 22833 28033 22845 28067
rect 22879 28064 22891 28067
rect 23198 28064 23204 28076
rect 22879 28036 23204 28064
rect 22879 28033 22891 28036
rect 22833 28027 22891 28033
rect 23198 28024 23204 28036
rect 23256 28024 23262 28076
rect 23293 28067 23351 28073
rect 23293 28033 23305 28067
rect 23339 28033 23351 28067
rect 23293 28027 23351 28033
rect 21818 27996 21824 28008
rect 21100 27968 21824 27996
rect 21818 27956 21824 27968
rect 21876 27956 21882 28008
rect 21910 27956 21916 28008
rect 21968 27956 21974 28008
rect 22281 27999 22339 28005
rect 22281 27996 22293 27999
rect 22066 27968 22293 27996
rect 21453 27931 21511 27937
rect 21008 27900 21312 27928
rect 21284 27872 21312 27900
rect 21453 27897 21465 27931
rect 21499 27928 21511 27931
rect 22066 27928 22094 27968
rect 22281 27965 22293 27968
rect 22327 27965 22339 27999
rect 22281 27959 22339 27965
rect 22741 27999 22799 28005
rect 22741 27965 22753 27999
rect 22787 27996 22799 27999
rect 22922 27996 22928 28008
rect 22787 27968 22928 27996
rect 22787 27965 22799 27968
rect 22741 27959 22799 27965
rect 22922 27956 22928 27968
rect 22980 27956 22986 28008
rect 23308 27996 23336 28027
rect 23382 28024 23388 28076
rect 23440 28024 23446 28076
rect 23477 28067 23535 28073
rect 23477 28033 23489 28067
rect 23523 28064 23535 28067
rect 23566 28064 23572 28076
rect 23523 28036 23572 28064
rect 23523 28033 23535 28036
rect 23477 28027 23535 28033
rect 23566 28024 23572 28036
rect 23624 28024 23630 28076
rect 23676 28073 23704 28104
rect 24688 28076 24716 28104
rect 31956 28104 34652 28132
rect 23661 28067 23719 28073
rect 23661 28033 23673 28067
rect 23707 28033 23719 28067
rect 23661 28027 23719 28033
rect 23750 28024 23756 28076
rect 23808 28024 23814 28076
rect 24026 28024 24032 28076
rect 24084 28064 24090 28076
rect 24121 28067 24179 28073
rect 24121 28064 24133 28067
rect 24084 28036 24133 28064
rect 24084 28024 24090 28036
rect 24121 28033 24133 28036
rect 24167 28033 24179 28067
rect 24121 28027 24179 28033
rect 24394 28024 24400 28076
rect 24452 28024 24458 28076
rect 24670 28024 24676 28076
rect 24728 28024 24734 28076
rect 31956 28073 31984 28104
rect 31941 28067 31999 28073
rect 31941 28033 31953 28067
rect 31987 28033 31999 28067
rect 32493 28067 32551 28073
rect 32493 28064 32505 28067
rect 31941 28027 31999 28033
rect 32232 28036 32505 28064
rect 23308 27968 23428 27996
rect 21499 27900 22094 27928
rect 21499 27897 21511 27900
rect 21453 27891 21511 27897
rect 20588 27832 20760 27860
rect 20588 27820 20594 27832
rect 21266 27820 21272 27872
rect 21324 27820 21330 27872
rect 22278 27820 22284 27872
rect 22336 27860 22342 27872
rect 23400 27860 23428 27968
rect 24029 27931 24087 27937
rect 24029 27897 24041 27931
rect 24075 27928 24087 27931
rect 24412 27928 24440 28024
rect 30190 27956 30196 28008
rect 30248 27996 30254 28008
rect 32232 27996 32260 28036
rect 32493 28033 32505 28036
rect 32539 28064 32551 28067
rect 34146 28064 34152 28076
rect 32539 28036 34152 28064
rect 32539 28033 32551 28036
rect 32493 28027 32551 28033
rect 34146 28024 34152 28036
rect 34204 28024 34210 28076
rect 34241 28067 34299 28073
rect 34241 28033 34253 28067
rect 34287 28064 34299 28067
rect 34514 28064 34520 28076
rect 34287 28036 34520 28064
rect 34287 28033 34299 28036
rect 34241 28027 34299 28033
rect 34514 28024 34520 28036
rect 34572 28024 34578 28076
rect 34624 28064 34652 28104
rect 34977 28067 35035 28073
rect 34977 28064 34989 28067
rect 34624 28036 34989 28064
rect 34977 28033 34989 28036
rect 35023 28033 35035 28067
rect 37292 28064 37320 28160
rect 37369 28067 37427 28073
rect 37369 28064 37381 28067
rect 37292 28036 37381 28064
rect 34977 28027 35035 28033
rect 37369 28033 37381 28036
rect 37415 28033 37427 28067
rect 37369 28027 37427 28033
rect 30248 27968 32260 27996
rect 32401 27999 32459 28005
rect 30248 27956 30254 27968
rect 32401 27965 32413 27999
rect 32447 27996 32459 27999
rect 33134 27996 33140 28008
rect 32447 27968 33140 27996
rect 32447 27965 32459 27968
rect 32401 27959 32459 27965
rect 33134 27956 33140 27968
rect 33192 27996 33198 28008
rect 33870 27996 33876 28008
rect 33192 27968 33876 27996
rect 33192 27956 33198 27968
rect 33870 27956 33876 27968
rect 33928 27956 33934 28008
rect 24075 27900 24440 27928
rect 24075 27897 24087 27900
rect 24029 27891 24087 27897
rect 22336 27832 23428 27860
rect 22336 27820 22342 27832
rect 24210 27820 24216 27872
rect 24268 27820 24274 27872
rect 24486 27820 24492 27872
rect 24544 27820 24550 27872
rect 26510 27820 26516 27872
rect 26568 27860 26574 27872
rect 28258 27860 28264 27872
rect 26568 27832 28264 27860
rect 26568 27820 26574 27832
rect 28258 27820 28264 27832
rect 28316 27820 28322 27872
rect 28810 27820 28816 27872
rect 28868 27860 28874 27872
rect 29730 27860 29736 27872
rect 28868 27832 29736 27860
rect 28868 27820 28874 27832
rect 29730 27820 29736 27832
rect 29788 27820 29794 27872
rect 37550 27820 37556 27872
rect 37608 27820 37614 27872
rect 1104 27770 38272 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38272 27770
rect 1104 27696 38272 27718
rect 4614 27616 4620 27668
rect 4672 27616 4678 27668
rect 8294 27616 8300 27668
rect 8352 27616 8358 27668
rect 9490 27616 9496 27668
rect 9548 27616 9554 27668
rect 9674 27616 9680 27668
rect 9732 27656 9738 27668
rect 9732 27628 14596 27656
rect 9732 27616 9738 27628
rect 9508 27588 9536 27616
rect 8496 27560 9536 27588
rect 4801 27455 4859 27461
rect 4801 27421 4813 27455
rect 4847 27452 4859 27455
rect 6362 27452 6368 27464
rect 4847 27424 6368 27452
rect 4847 27421 4859 27424
rect 4801 27415 4859 27421
rect 6362 27412 6368 27424
rect 6420 27412 6426 27464
rect 6914 27412 6920 27464
rect 6972 27452 6978 27464
rect 8496 27461 8524 27560
rect 9582 27548 9588 27600
rect 9640 27548 9646 27600
rect 14090 27548 14096 27600
rect 14148 27548 14154 27600
rect 14568 27588 14596 27628
rect 14642 27616 14648 27668
rect 14700 27616 14706 27668
rect 14752 27628 15976 27656
rect 14752 27588 14780 27628
rect 14568 27560 14780 27588
rect 15948 27588 15976 27628
rect 16022 27616 16028 27668
rect 16080 27616 16086 27668
rect 20438 27656 20444 27668
rect 16132 27628 20444 27656
rect 16132 27588 16160 27628
rect 20438 27616 20444 27628
rect 20496 27656 20502 27668
rect 23382 27656 23388 27668
rect 20496 27628 23388 27656
rect 20496 27616 20502 27628
rect 17126 27588 17132 27600
rect 15948 27560 16160 27588
rect 16868 27560 17132 27588
rect 9600 27520 9628 27548
rect 9508 27492 9628 27520
rect 9508 27461 9536 27492
rect 11974 27480 11980 27532
rect 12032 27520 12038 27532
rect 12069 27523 12127 27529
rect 12069 27520 12081 27523
rect 12032 27492 12081 27520
rect 12032 27480 12038 27492
rect 12069 27489 12081 27492
rect 12115 27489 12127 27523
rect 12069 27483 12127 27489
rect 12253 27523 12311 27529
rect 12253 27489 12265 27523
rect 12299 27520 12311 27523
rect 13081 27523 13139 27529
rect 12299 27492 12434 27520
rect 12299 27489 12311 27492
rect 12253 27483 12311 27489
rect 8481 27455 8539 27461
rect 6972 27424 7604 27452
rect 6972 27412 6978 27424
rect 7576 27328 7604 27424
rect 8481 27421 8493 27455
rect 8527 27421 8539 27455
rect 8481 27415 8539 27421
rect 9493 27455 9551 27461
rect 9493 27421 9505 27455
rect 9539 27421 9551 27455
rect 9493 27415 9551 27421
rect 9585 27455 9643 27461
rect 9585 27421 9597 27455
rect 9631 27452 9643 27455
rect 9769 27455 9827 27461
rect 9769 27452 9781 27455
rect 9631 27424 9781 27452
rect 9631 27421 9643 27424
rect 9585 27415 9643 27421
rect 9769 27421 9781 27424
rect 9815 27421 9827 27455
rect 9769 27415 9827 27421
rect 11054 27412 11060 27464
rect 11112 27452 11118 27464
rect 11112 27424 11178 27452
rect 11112 27412 11118 27424
rect 10042 27344 10048 27396
rect 10100 27344 10106 27396
rect 12406 27384 12434 27492
rect 13081 27489 13093 27523
rect 13127 27520 13139 27523
rect 13722 27520 13728 27532
rect 13127 27492 13728 27520
rect 13127 27489 13139 27492
rect 13081 27483 13139 27489
rect 13722 27480 13728 27492
rect 13780 27480 13786 27532
rect 13170 27412 13176 27464
rect 13228 27452 13234 27464
rect 13265 27455 13323 27461
rect 13265 27452 13277 27455
rect 13228 27424 13277 27452
rect 13228 27412 13234 27424
rect 13265 27421 13277 27424
rect 13311 27452 13323 27455
rect 13538 27452 13544 27464
rect 13311 27424 13544 27452
rect 13311 27421 13323 27424
rect 13265 27415 13323 27421
rect 13538 27412 13544 27424
rect 13596 27412 13602 27464
rect 13814 27412 13820 27464
rect 13872 27412 13878 27464
rect 15562 27412 15568 27464
rect 15620 27412 15626 27464
rect 15657 27455 15715 27461
rect 15657 27421 15669 27455
rect 15703 27421 15715 27455
rect 15657 27415 15715 27421
rect 15841 27455 15899 27461
rect 15841 27421 15853 27455
rect 15887 27452 15899 27455
rect 16114 27452 16120 27464
rect 15887 27424 16120 27452
rect 15887 27421 15899 27424
rect 15841 27415 15899 27421
rect 12526 27384 12532 27396
rect 11532 27356 12020 27384
rect 12406 27356 12532 27384
rect 6822 27276 6828 27328
rect 6880 27276 6886 27328
rect 7558 27276 7564 27328
rect 7616 27276 7622 27328
rect 11532 27325 11560 27356
rect 11517 27319 11575 27325
rect 11517 27285 11529 27319
rect 11563 27285 11575 27319
rect 11517 27279 11575 27285
rect 11606 27276 11612 27328
rect 11664 27276 11670 27328
rect 11992 27325 12020 27356
rect 12526 27344 12532 27356
rect 12584 27344 12590 27396
rect 13832 27384 13860 27412
rect 14458 27384 14464 27396
rect 13832 27356 14464 27384
rect 14458 27344 14464 27356
rect 14516 27344 14522 27396
rect 15672 27384 15700 27415
rect 16114 27412 16120 27424
rect 16172 27412 16178 27464
rect 16574 27412 16580 27464
rect 16632 27412 16638 27464
rect 16666 27412 16672 27464
rect 16724 27412 16730 27464
rect 16758 27412 16764 27464
rect 16816 27412 16822 27464
rect 16868 27452 16896 27560
rect 17126 27548 17132 27560
rect 17184 27548 17190 27600
rect 17586 27588 17592 27600
rect 17236 27560 17592 27588
rect 17236 27520 17264 27560
rect 17586 27548 17592 27560
rect 17644 27548 17650 27600
rect 17678 27548 17684 27600
rect 17736 27588 17742 27600
rect 18966 27588 18972 27600
rect 17736 27560 18972 27588
rect 17736 27548 17742 27560
rect 18966 27548 18972 27560
rect 19024 27548 19030 27600
rect 20162 27548 20168 27600
rect 20220 27588 20226 27600
rect 20622 27588 20628 27600
rect 20220 27560 20628 27588
rect 20220 27548 20226 27560
rect 20622 27548 20628 27560
rect 20680 27548 20686 27600
rect 17139 27492 17264 27520
rect 17139 27461 17167 27492
rect 17862 27480 17868 27532
rect 17920 27480 17926 27532
rect 18046 27480 18052 27532
rect 18104 27520 18110 27532
rect 21266 27520 21272 27532
rect 18104 27492 21272 27520
rect 18104 27480 18110 27492
rect 17402 27461 17408 27464
rect 16945 27455 17003 27461
rect 16945 27452 16957 27455
rect 16868 27424 16957 27452
rect 16945 27421 16957 27424
rect 16991 27421 17003 27455
rect 16945 27415 17003 27421
rect 17134 27455 17192 27461
rect 17134 27421 17146 27455
rect 17180 27421 17192 27455
rect 17134 27415 17192 27421
rect 17393 27455 17408 27461
rect 17393 27421 17405 27455
rect 17393 27415 17408 27421
rect 17402 27412 17408 27415
rect 17460 27412 17466 27464
rect 17494 27412 17500 27464
rect 17552 27452 17558 27464
rect 17589 27455 17647 27461
rect 17589 27452 17601 27455
rect 17552 27424 17601 27452
rect 17552 27412 17558 27424
rect 17589 27421 17601 27424
rect 17635 27421 17647 27455
rect 17589 27415 17647 27421
rect 17678 27412 17684 27464
rect 17736 27412 17742 27464
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27452 17831 27455
rect 17880 27452 17908 27480
rect 17819 27424 17908 27452
rect 17819 27421 17831 27424
rect 17773 27415 17831 27421
rect 18138 27412 18144 27464
rect 18196 27412 18202 27464
rect 18432 27461 18460 27492
rect 21266 27480 21272 27492
rect 21324 27520 21330 27532
rect 21726 27520 21732 27532
rect 21324 27492 21732 27520
rect 21324 27480 21330 27492
rect 21726 27480 21732 27492
rect 21784 27480 21790 27532
rect 18325 27455 18383 27461
rect 18325 27421 18337 27455
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 18417 27455 18475 27461
rect 18417 27421 18429 27455
rect 18463 27421 18475 27455
rect 18417 27415 18475 27421
rect 16592 27384 16620 27412
rect 15672 27356 16620 27384
rect 17037 27387 17095 27393
rect 17037 27353 17049 27387
rect 17083 27353 17095 27387
rect 17037 27347 17095 27353
rect 18049 27387 18107 27393
rect 18049 27353 18061 27387
rect 18095 27384 18107 27387
rect 18340 27384 18368 27415
rect 18598 27412 18604 27464
rect 18656 27412 18662 27464
rect 19334 27412 19340 27464
rect 19392 27452 19398 27464
rect 22940 27461 22968 27628
rect 23382 27616 23388 27628
rect 23440 27616 23446 27668
rect 23753 27659 23811 27665
rect 23753 27625 23765 27659
rect 23799 27656 23811 27659
rect 24210 27656 24216 27668
rect 23799 27628 24216 27656
rect 23799 27625 23811 27628
rect 23753 27619 23811 27625
rect 24210 27616 24216 27628
rect 24268 27616 24274 27668
rect 24394 27656 24400 27668
rect 24320 27628 24400 27656
rect 23566 27588 23572 27600
rect 23032 27560 23572 27588
rect 22925 27455 22983 27461
rect 19392 27424 22876 27452
rect 19392 27412 19398 27424
rect 18095 27356 18368 27384
rect 18095 27353 18107 27356
rect 18049 27347 18107 27353
rect 11977 27319 12035 27325
rect 11977 27285 11989 27319
rect 12023 27316 12035 27319
rect 12342 27316 12348 27328
rect 12023 27288 12348 27316
rect 12023 27285 12035 27288
rect 11977 27279 12035 27285
rect 12342 27276 12348 27288
rect 12400 27276 12406 27328
rect 14274 27276 14280 27328
rect 14332 27276 14338 27328
rect 14366 27276 14372 27328
rect 14424 27316 14430 27328
rect 14550 27316 14556 27328
rect 14424 27288 14556 27316
rect 14424 27276 14430 27288
rect 14550 27276 14556 27288
rect 14608 27276 14614 27328
rect 15562 27276 15568 27328
rect 15620 27316 15626 27328
rect 16850 27316 16856 27328
rect 15620 27288 16856 27316
rect 15620 27276 15626 27288
rect 16850 27276 16856 27288
rect 16908 27316 16914 27328
rect 17052 27316 17080 27347
rect 18506 27344 18512 27396
rect 18564 27344 18570 27396
rect 19426 27384 19432 27396
rect 18708 27356 19432 27384
rect 16908 27288 17080 27316
rect 17313 27319 17371 27325
rect 16908 27276 16914 27288
rect 17313 27285 17325 27319
rect 17359 27316 17371 27319
rect 17770 27316 17776 27328
rect 17359 27288 17776 27316
rect 17359 27285 17371 27288
rect 17313 27279 17371 27285
rect 17770 27276 17776 27288
rect 17828 27276 17834 27328
rect 18414 27276 18420 27328
rect 18472 27316 18478 27328
rect 18708 27316 18736 27356
rect 19426 27344 19432 27356
rect 19484 27344 19490 27396
rect 19886 27344 19892 27396
rect 19944 27384 19950 27396
rect 21082 27384 21088 27396
rect 19944 27356 21088 27384
rect 19944 27344 19950 27356
rect 21082 27344 21088 27356
rect 21140 27384 21146 27396
rect 21450 27384 21456 27396
rect 21140 27356 21456 27384
rect 21140 27344 21146 27356
rect 21450 27344 21456 27356
rect 21508 27344 21514 27396
rect 22741 27387 22799 27393
rect 22741 27384 22753 27387
rect 22066 27356 22753 27384
rect 18472 27288 18736 27316
rect 18472 27276 18478 27288
rect 18782 27276 18788 27328
rect 18840 27276 18846 27328
rect 20162 27276 20168 27328
rect 20220 27316 20226 27328
rect 22066 27316 22094 27356
rect 22741 27353 22753 27356
rect 22787 27353 22799 27387
rect 22848 27384 22876 27424
rect 22925 27421 22937 27455
rect 22971 27421 22983 27455
rect 22925 27415 22983 27421
rect 23032 27384 23060 27560
rect 23566 27548 23572 27560
rect 23624 27548 23630 27600
rect 24320 27520 24348 27628
rect 24394 27616 24400 27628
rect 24452 27656 24458 27668
rect 26694 27656 26700 27668
rect 24452 27628 26700 27656
rect 24452 27616 24458 27628
rect 26694 27616 26700 27628
rect 26752 27616 26758 27668
rect 27614 27616 27620 27668
rect 27672 27656 27678 27668
rect 34606 27656 34612 27668
rect 27672 27628 28396 27656
rect 27672 27616 27678 27628
rect 28368 27600 28396 27628
rect 33704 27628 34612 27656
rect 25498 27548 25504 27600
rect 25556 27548 25562 27600
rect 28350 27548 28356 27600
rect 28408 27548 28414 27600
rect 30300 27560 30788 27588
rect 23216 27492 24348 27520
rect 23216 27461 23244 27492
rect 23201 27455 23259 27461
rect 23201 27421 23213 27455
rect 23247 27421 23259 27455
rect 23201 27415 23259 27421
rect 23477 27455 23535 27461
rect 23477 27421 23489 27455
rect 23523 27421 23535 27455
rect 23477 27415 23535 27421
rect 22848 27356 23060 27384
rect 23109 27387 23167 27393
rect 22741 27347 22799 27353
rect 23109 27353 23121 27387
rect 23155 27384 23167 27387
rect 23385 27387 23443 27393
rect 23385 27384 23397 27387
rect 23155 27356 23397 27384
rect 23155 27353 23167 27356
rect 23109 27347 23167 27353
rect 23385 27353 23397 27356
rect 23431 27353 23443 27387
rect 23385 27347 23443 27353
rect 20220 27288 22094 27316
rect 20220 27276 20226 27288
rect 22186 27276 22192 27328
rect 22244 27316 22250 27328
rect 23492 27316 23520 27415
rect 23566 27412 23572 27464
rect 23624 27412 23630 27464
rect 25516 27461 25544 27548
rect 29086 27520 29092 27532
rect 27908 27492 29092 27520
rect 27908 27461 27936 27492
rect 29086 27480 29092 27492
rect 29144 27520 29150 27532
rect 29638 27520 29644 27532
rect 29144 27492 29644 27520
rect 29144 27480 29150 27492
rect 29638 27480 29644 27492
rect 29696 27480 29702 27532
rect 25501 27455 25559 27461
rect 25501 27421 25513 27455
rect 25547 27421 25559 27455
rect 25501 27415 25559 27421
rect 25593 27455 25651 27461
rect 25593 27421 25605 27455
rect 25639 27452 25651 27455
rect 25777 27455 25835 27461
rect 25777 27452 25789 27455
rect 25639 27424 25789 27452
rect 25639 27421 25651 27424
rect 25593 27415 25651 27421
rect 25777 27421 25789 27424
rect 25823 27421 25835 27455
rect 25777 27415 25835 27421
rect 27893 27455 27951 27461
rect 27893 27421 27905 27455
rect 27939 27421 27951 27455
rect 27893 27415 27951 27421
rect 28166 27412 28172 27464
rect 28224 27412 28230 27464
rect 29178 27452 29184 27464
rect 28276 27424 29184 27452
rect 26050 27344 26056 27396
rect 26108 27344 26114 27396
rect 27430 27384 27436 27396
rect 27278 27356 27436 27384
rect 27430 27344 27436 27356
rect 27488 27384 27494 27396
rect 28276 27384 28304 27424
rect 29178 27412 29184 27424
rect 29236 27412 29242 27464
rect 29549 27455 29607 27461
rect 29549 27421 29561 27455
rect 29595 27452 29607 27455
rect 29656 27452 29684 27480
rect 29595 27424 29684 27452
rect 29595 27421 29607 27424
rect 29549 27415 29607 27421
rect 30006 27412 30012 27464
rect 30064 27412 30070 27464
rect 30300 27384 30328 27560
rect 30374 27412 30380 27464
rect 30432 27412 30438 27464
rect 30470 27455 30528 27461
rect 30470 27421 30482 27455
rect 30516 27421 30528 27455
rect 30470 27415 30528 27421
rect 30484 27384 30512 27415
rect 30650 27412 30656 27464
rect 30708 27412 30714 27464
rect 30760 27393 30788 27560
rect 30926 27461 30932 27464
rect 30883 27455 30932 27461
rect 30883 27421 30895 27455
rect 30929 27421 30932 27455
rect 30883 27415 30932 27421
rect 30926 27412 30932 27415
rect 30984 27412 30990 27464
rect 33704 27461 33732 27628
rect 34606 27616 34612 27628
rect 34664 27616 34670 27668
rect 33778 27548 33784 27600
rect 33836 27548 33842 27600
rect 34330 27548 34336 27600
rect 34388 27548 34394 27600
rect 33689 27455 33747 27461
rect 33689 27421 33701 27455
rect 33735 27421 33747 27455
rect 33689 27415 33747 27421
rect 33965 27455 34023 27461
rect 33965 27421 33977 27455
rect 34011 27452 34023 27455
rect 34348 27452 34376 27548
rect 34011 27424 34376 27452
rect 34011 27421 34023 27424
rect 33965 27415 34023 27421
rect 27488 27356 28304 27384
rect 28966 27356 30328 27384
rect 30392 27356 30512 27384
rect 30745 27387 30803 27393
rect 27488 27344 27494 27356
rect 22244 27288 23520 27316
rect 22244 27276 22250 27288
rect 26418 27276 26424 27328
rect 26476 27316 26482 27328
rect 27525 27319 27583 27325
rect 27525 27316 27537 27319
rect 26476 27288 27537 27316
rect 26476 27276 26482 27288
rect 27525 27285 27537 27288
rect 27571 27285 27583 27319
rect 27525 27279 27583 27285
rect 27798 27276 27804 27328
rect 27856 27276 27862 27328
rect 27890 27276 27896 27328
rect 27948 27316 27954 27328
rect 27985 27319 28043 27325
rect 27985 27316 27997 27319
rect 27948 27288 27997 27316
rect 27948 27276 27954 27288
rect 27985 27285 27997 27288
rect 28031 27285 28043 27319
rect 27985 27279 28043 27285
rect 28258 27276 28264 27328
rect 28316 27316 28322 27328
rect 28966 27316 28994 27356
rect 30392 27328 30420 27356
rect 30745 27353 30757 27387
rect 30791 27384 30803 27387
rect 32674 27384 32680 27396
rect 30791 27356 32680 27384
rect 30791 27353 30803 27356
rect 30745 27347 30803 27353
rect 32674 27344 32680 27356
rect 32732 27344 32738 27396
rect 28316 27288 28994 27316
rect 28316 27276 28322 27288
rect 29638 27276 29644 27328
rect 29696 27276 29702 27328
rect 29822 27276 29828 27328
rect 29880 27276 29886 27328
rect 30374 27276 30380 27328
rect 30432 27276 30438 27328
rect 31021 27319 31079 27325
rect 31021 27285 31033 27319
rect 31067 27316 31079 27319
rect 31754 27316 31760 27328
rect 31067 27288 31760 27316
rect 31067 27285 31079 27288
rect 31021 27279 31079 27285
rect 31754 27276 31760 27288
rect 31812 27276 31818 27328
rect 33594 27276 33600 27328
rect 33652 27276 33658 27328
rect 1104 27226 38272 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38272 27226
rect 1104 27152 38272 27174
rect 6822 27072 6828 27124
rect 6880 27072 6886 27124
rect 10042 27072 10048 27124
rect 10100 27112 10106 27124
rect 10229 27115 10287 27121
rect 10229 27112 10241 27115
rect 10100 27084 10241 27112
rect 10100 27072 10106 27084
rect 10229 27081 10241 27084
rect 10275 27081 10287 27115
rect 10229 27075 10287 27081
rect 11606 27072 11612 27124
rect 11664 27072 11670 27124
rect 12158 27072 12164 27124
rect 12216 27112 12222 27124
rect 16298 27112 16304 27124
rect 12216 27084 12802 27112
rect 12216 27072 12222 27084
rect 6840 27044 6868 27072
rect 6656 27016 6868 27044
rect 6656 26985 6684 27016
rect 7190 27004 7196 27056
rect 7248 27044 7254 27056
rect 7374 27044 7380 27056
rect 7248 27016 7380 27044
rect 7248 27004 7254 27016
rect 7374 27004 7380 27016
rect 7432 27004 7438 27056
rect 6641 26979 6699 26985
rect 6641 26945 6653 26979
rect 6687 26945 6699 26979
rect 6641 26939 6699 26945
rect 10413 26979 10471 26985
rect 10413 26945 10425 26979
rect 10459 26976 10471 26979
rect 11624 26976 11652 27072
rect 11882 27004 11888 27056
rect 11940 27044 11946 27056
rect 12529 27047 12587 27053
rect 12529 27044 12541 27047
rect 11940 27016 12541 27044
rect 11940 27004 11946 27016
rect 12529 27013 12541 27016
rect 12575 27013 12587 27047
rect 12529 27007 12587 27013
rect 12774 26988 12802 27084
rect 13924 27084 16304 27112
rect 10459 26948 11652 26976
rect 10459 26945 10471 26948
rect 10413 26939 10471 26945
rect 12250 26936 12256 26988
rect 12308 26936 12314 26988
rect 12342 26936 12348 26988
rect 12400 26976 12406 26988
rect 12774 26985 12808 26988
rect 12621 26979 12679 26985
rect 12400 26948 12445 26976
rect 12400 26936 12406 26948
rect 12621 26945 12633 26979
rect 12667 26945 12679 26979
rect 12621 26939 12679 26945
rect 12759 26979 12808 26985
rect 12759 26945 12771 26979
rect 12805 26945 12808 26979
rect 12759 26939 12808 26945
rect 6914 26868 6920 26920
rect 6972 26868 6978 26920
rect 7466 26868 7472 26920
rect 7524 26908 7530 26920
rect 7524 26880 8340 26908
rect 7524 26868 7530 26880
rect 8312 26840 8340 26880
rect 8386 26868 8392 26920
rect 8444 26908 8450 26920
rect 12636 26908 12664 26939
rect 12802 26936 12808 26939
rect 12860 26976 12866 26988
rect 13924 26976 13952 27084
rect 16298 27072 16304 27084
rect 16356 27072 16362 27124
rect 16666 27072 16672 27124
rect 16724 27072 16730 27124
rect 16942 27072 16948 27124
rect 17000 27072 17006 27124
rect 18049 27115 18107 27121
rect 17236 27084 18000 27112
rect 13998 27004 14004 27056
rect 14056 27004 14062 27056
rect 14366 27004 14372 27056
rect 14424 27044 14430 27056
rect 14642 27044 14648 27056
rect 14424 27016 14648 27044
rect 14424 27004 14430 27016
rect 14642 27004 14648 27016
rect 14700 27004 14706 27056
rect 15470 27004 15476 27056
rect 15528 27004 15534 27056
rect 17236 27044 17264 27084
rect 15580 27016 17264 27044
rect 12860 26948 13952 26976
rect 14016 26976 14044 27004
rect 14461 26979 14519 26985
rect 14461 26976 14473 26979
rect 14016 26948 14473 26976
rect 12860 26936 12866 26948
rect 14461 26945 14473 26948
rect 14507 26945 14519 26979
rect 14461 26939 14519 26945
rect 14734 26936 14740 26988
rect 14792 26936 14798 26988
rect 14921 26979 14979 26985
rect 14921 26945 14933 26979
rect 14967 26976 14979 26979
rect 15010 26976 15016 26988
rect 14967 26948 15016 26976
rect 14967 26945 14979 26948
rect 14921 26939 14979 26945
rect 15010 26936 15016 26948
rect 15068 26936 15074 26988
rect 15378 26936 15384 26988
rect 15436 26976 15442 26988
rect 15580 26976 15608 27016
rect 15436 26948 15608 26976
rect 15436 26936 15442 26948
rect 15654 26936 15660 26988
rect 15712 26936 15718 26988
rect 16390 26936 16396 26988
rect 16448 26976 16454 26988
rect 16758 26976 16764 26988
rect 16448 26948 16764 26976
rect 16448 26936 16454 26948
rect 16758 26936 16764 26948
rect 16816 26936 16822 26988
rect 16853 26979 16911 26985
rect 16853 26945 16865 26979
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 8444 26880 14509 26908
rect 8444 26868 8450 26880
rect 9858 26840 9864 26852
rect 8312 26812 9864 26840
rect 9858 26800 9864 26812
rect 9916 26840 9922 26852
rect 12526 26840 12532 26852
rect 9916 26812 12532 26840
rect 9916 26800 9922 26812
rect 12526 26800 12532 26812
rect 12584 26840 12590 26852
rect 14182 26840 14188 26852
rect 12584 26812 14188 26840
rect 12584 26800 12590 26812
rect 14182 26800 14188 26812
rect 14240 26800 14246 26852
rect 5994 26732 6000 26784
rect 6052 26772 6058 26784
rect 7374 26772 7380 26784
rect 6052 26744 7380 26772
rect 6052 26732 6058 26744
rect 7374 26732 7380 26744
rect 7432 26732 7438 26784
rect 12894 26732 12900 26784
rect 12952 26732 12958 26784
rect 14274 26732 14280 26784
rect 14332 26732 14338 26784
rect 14481 26772 14509 26880
rect 14642 26868 14648 26920
rect 14700 26868 14706 26920
rect 15470 26868 15476 26920
rect 15528 26908 15534 26920
rect 16408 26908 16436 26936
rect 15528 26880 16436 26908
rect 15528 26868 15534 26880
rect 14553 26843 14611 26849
rect 14553 26809 14565 26843
rect 14599 26840 14611 26843
rect 15102 26840 15108 26852
rect 14599 26812 15108 26840
rect 14599 26809 14611 26812
rect 14553 26803 14611 26809
rect 15102 26800 15108 26812
rect 15160 26800 15166 26852
rect 16868 26840 16896 26939
rect 17034 26936 17040 26988
rect 17092 26976 17098 26988
rect 17218 26976 17224 26988
rect 17092 26948 17224 26976
rect 17092 26936 17098 26948
rect 17218 26936 17224 26948
rect 17276 26936 17282 26988
rect 17678 26936 17684 26988
rect 17736 26936 17742 26988
rect 17770 26936 17776 26988
rect 17828 26936 17834 26988
rect 17972 26976 18000 27084
rect 18049 27081 18061 27115
rect 18095 27112 18107 27115
rect 18506 27112 18512 27124
rect 18095 27084 18512 27112
rect 18095 27081 18107 27084
rect 18049 27075 18107 27081
rect 18506 27072 18512 27084
rect 18564 27072 18570 27124
rect 18598 27072 18604 27124
rect 18656 27112 18662 27124
rect 18785 27115 18843 27121
rect 18785 27112 18797 27115
rect 18656 27084 18797 27112
rect 18656 27072 18662 27084
rect 18785 27081 18797 27084
rect 18831 27081 18843 27115
rect 18785 27075 18843 27081
rect 18966 27072 18972 27124
rect 19024 27072 19030 27124
rect 22186 27072 22192 27124
rect 22244 27072 22250 27124
rect 24762 27112 24768 27124
rect 22388 27084 24768 27112
rect 18984 27044 19012 27072
rect 18984 27016 19196 27044
rect 17972 26948 18920 26976
rect 16942 26868 16948 26920
rect 17000 26908 17006 26920
rect 18506 26908 18512 26920
rect 17000 26880 18512 26908
rect 17000 26868 17006 26880
rect 18506 26868 18512 26880
rect 18564 26868 18570 26920
rect 18892 26908 18920 26948
rect 18966 26936 18972 26988
rect 19024 26936 19030 26988
rect 19168 26985 19196 27016
rect 19153 26979 19211 26985
rect 19153 26945 19165 26979
rect 19199 26945 19211 26979
rect 19153 26939 19211 26945
rect 19426 26936 19432 26988
rect 19484 26936 19490 26988
rect 22388 26985 22416 27084
rect 24762 27072 24768 27084
rect 24820 27072 24826 27124
rect 26050 27072 26056 27124
rect 26108 27112 26114 27124
rect 26973 27115 27031 27121
rect 26973 27112 26985 27115
rect 26108 27084 26985 27112
rect 26108 27072 26114 27084
rect 26973 27081 26985 27084
rect 27019 27081 27031 27115
rect 26973 27075 27031 27081
rect 27798 27072 27804 27124
rect 27856 27072 27862 27124
rect 28626 27072 28632 27124
rect 28684 27112 28690 27124
rect 28684 27084 28948 27112
rect 28684 27072 28690 27084
rect 22557 27047 22615 27053
rect 22557 27013 22569 27047
rect 22603 27044 22615 27047
rect 23474 27044 23480 27056
rect 22603 27016 23480 27044
rect 22603 27013 22615 27016
rect 22557 27007 22615 27013
rect 23474 27004 23480 27016
rect 23532 27004 23538 27056
rect 26329 27047 26387 27053
rect 26329 27013 26341 27047
rect 26375 27044 26387 27047
rect 27816 27044 27844 27072
rect 26375 27016 27384 27044
rect 26375 27013 26387 27016
rect 26329 27007 26387 27013
rect 22373 26979 22431 26985
rect 22373 26945 22385 26979
rect 22419 26945 22431 26979
rect 22373 26939 22431 26945
rect 22465 26979 22523 26985
rect 22465 26945 22477 26979
rect 22511 26945 22523 26979
rect 22465 26939 22523 26945
rect 19334 26908 19340 26920
rect 18892 26880 19340 26908
rect 19334 26868 19340 26880
rect 19392 26868 19398 26920
rect 19444 26908 19472 26936
rect 22480 26908 22508 26939
rect 22738 26936 22744 26988
rect 22796 26936 22802 26988
rect 24670 26936 24676 26988
rect 24728 26976 24734 26988
rect 25958 26976 25964 26988
rect 24728 26948 25964 26976
rect 24728 26936 24734 26948
rect 25958 26936 25964 26948
rect 26016 26936 26022 26988
rect 26418 26976 26424 26988
rect 26068 26948 26424 26976
rect 24762 26908 24768 26920
rect 19444 26880 24768 26908
rect 24762 26868 24768 26880
rect 24820 26908 24826 26920
rect 26068 26908 26096 26948
rect 26418 26936 26424 26948
rect 26476 26936 26482 26988
rect 27157 26979 27215 26985
rect 27157 26976 27169 26979
rect 26804 26948 27169 26976
rect 24820 26880 26096 26908
rect 26237 26911 26295 26917
rect 24820 26868 24826 26880
rect 26237 26877 26249 26911
rect 26283 26908 26295 26911
rect 26510 26908 26516 26920
rect 26283 26880 26516 26908
rect 26283 26877 26295 26880
rect 26237 26871 26295 26877
rect 26510 26868 26516 26880
rect 26568 26868 26574 26920
rect 17126 26840 17132 26852
rect 16868 26812 17132 26840
rect 17126 26800 17132 26812
rect 17184 26800 17190 26852
rect 17221 26843 17279 26849
rect 17221 26809 17233 26843
rect 17267 26840 17279 26843
rect 17310 26840 17316 26852
rect 17267 26812 17316 26840
rect 17267 26809 17279 26812
rect 17221 26803 17279 26809
rect 17310 26800 17316 26812
rect 17368 26840 17374 26852
rect 26050 26840 26056 26852
rect 17368 26812 26056 26840
rect 17368 26800 17374 26812
rect 26050 26800 26056 26812
rect 26108 26800 26114 26852
rect 26804 26849 26832 26948
rect 27157 26945 27169 26948
rect 27203 26945 27215 26979
rect 27157 26939 27215 26945
rect 27356 26920 27384 27016
rect 27540 27016 27844 27044
rect 27540 26985 27568 27016
rect 27525 26979 27583 26985
rect 27525 26945 27537 26979
rect 27571 26945 27583 26979
rect 27525 26939 27583 26945
rect 27338 26868 27344 26920
rect 27396 26868 27402 26920
rect 27801 26911 27859 26917
rect 27801 26877 27813 26911
rect 27847 26908 27859 26911
rect 27890 26908 27896 26920
rect 27847 26880 27896 26908
rect 27847 26877 27859 26880
rect 27801 26871 27859 26877
rect 27890 26868 27896 26880
rect 27948 26868 27954 26920
rect 28920 26908 28948 27084
rect 29638 27072 29644 27124
rect 29696 27072 29702 27124
rect 29822 27112 29828 27124
rect 29748 27084 29828 27112
rect 29656 27044 29684 27072
rect 29748 27053 29776 27084
rect 29822 27072 29828 27084
rect 29880 27072 29886 27124
rect 31570 27112 31576 27124
rect 31312 27084 31576 27112
rect 29472 27016 29684 27044
rect 29733 27047 29791 27053
rect 29472 26985 29500 27016
rect 29733 27013 29745 27047
rect 29779 27013 29791 27047
rect 29733 27007 29791 27013
rect 29457 26979 29515 26985
rect 29457 26945 29469 26979
rect 29503 26945 29515 26979
rect 31312 26976 31340 27084
rect 31570 27072 31576 27084
rect 31628 27112 31634 27124
rect 34054 27112 34060 27124
rect 31628 27084 34060 27112
rect 31628 27072 31634 27084
rect 34054 27072 34060 27084
rect 34112 27112 34118 27124
rect 34112 27084 34836 27112
rect 34112 27072 34118 27084
rect 33594 27044 33600 27056
rect 33428 27016 33600 27044
rect 30866 26962 31340 26976
rect 29457 26939 29515 26945
rect 30852 26948 31340 26962
rect 29730 26908 29736 26920
rect 28920 26880 29736 26908
rect 29730 26868 29736 26880
rect 29788 26908 29794 26920
rect 30852 26908 30880 26948
rect 31662 26936 31668 26988
rect 31720 26936 31726 26988
rect 33134 26936 33140 26988
rect 33192 26936 33198 26988
rect 33428 26985 33456 27016
rect 33594 27004 33600 27016
rect 33652 27004 33658 27056
rect 33413 26979 33471 26985
rect 33413 26945 33425 26979
rect 33459 26945 33471 26979
rect 34808 26976 34836 27084
rect 35986 26976 35992 26988
rect 34808 26962 35992 26976
rect 34822 26948 35992 26962
rect 33413 26939 33471 26945
rect 35986 26936 35992 26948
rect 36044 26936 36050 26988
rect 33689 26911 33747 26917
rect 33689 26908 33701 26911
rect 29788 26880 30880 26908
rect 33336 26880 33701 26908
rect 29788 26868 29794 26880
rect 26789 26843 26847 26849
rect 26789 26809 26801 26843
rect 26835 26809 26847 26843
rect 26789 26803 26847 26809
rect 28994 26800 29000 26852
rect 29052 26840 29058 26852
rect 33336 26849 33364 26880
rect 33689 26877 33701 26880
rect 33735 26877 33747 26911
rect 33689 26871 33747 26877
rect 33778 26868 33784 26920
rect 33836 26908 33842 26920
rect 35437 26911 35495 26917
rect 35437 26908 35449 26911
rect 33836 26880 35449 26908
rect 33836 26868 33842 26880
rect 35437 26877 35449 26880
rect 35483 26877 35495 26911
rect 35437 26871 35495 26877
rect 33321 26843 33379 26849
rect 29052 26812 29592 26840
rect 29052 26800 29058 26812
rect 15562 26772 15568 26784
rect 14481 26744 15568 26772
rect 15562 26732 15568 26744
rect 15620 26732 15626 26784
rect 16942 26732 16948 26784
rect 17000 26772 17006 26784
rect 17494 26772 17500 26784
rect 17000 26744 17500 26772
rect 17000 26732 17006 26744
rect 17494 26732 17500 26744
rect 17552 26732 17558 26784
rect 17678 26732 17684 26784
rect 17736 26732 17742 26784
rect 18874 26732 18880 26784
rect 18932 26772 18938 26784
rect 18969 26775 19027 26781
rect 18969 26772 18981 26775
rect 18932 26744 18981 26772
rect 18932 26732 18938 26744
rect 18969 26741 18981 26744
rect 19015 26741 19027 26775
rect 18969 26735 19027 26741
rect 19334 26732 19340 26784
rect 19392 26772 19398 26784
rect 19978 26772 19984 26784
rect 19392 26744 19984 26772
rect 19392 26732 19398 26744
rect 19978 26732 19984 26744
rect 20036 26732 20042 26784
rect 22554 26732 22560 26784
rect 22612 26772 22618 26784
rect 25866 26772 25872 26784
rect 22612 26744 25872 26772
rect 22612 26732 22618 26744
rect 25866 26732 25872 26744
rect 25924 26732 25930 26784
rect 28258 26732 28264 26784
rect 28316 26772 28322 26784
rect 29273 26775 29331 26781
rect 29273 26772 29285 26775
rect 28316 26744 29285 26772
rect 28316 26732 28322 26744
rect 29273 26741 29285 26744
rect 29319 26741 29331 26775
rect 29564 26772 29592 26812
rect 33321 26809 33333 26843
rect 33367 26809 33379 26843
rect 33321 26803 33379 26809
rect 30374 26772 30380 26784
rect 29564 26744 30380 26772
rect 29273 26735 29331 26741
rect 30374 26732 30380 26744
rect 30432 26772 30438 26784
rect 31205 26775 31263 26781
rect 31205 26772 31217 26775
rect 30432 26744 31217 26772
rect 30432 26732 30438 26744
rect 31205 26741 31217 26744
rect 31251 26741 31263 26775
rect 31205 26735 31263 26741
rect 31386 26732 31392 26784
rect 31444 26772 31450 26784
rect 31481 26775 31539 26781
rect 31481 26772 31493 26775
rect 31444 26744 31493 26772
rect 31444 26732 31450 26744
rect 31481 26741 31493 26744
rect 31527 26741 31539 26775
rect 31481 26735 31539 26741
rect 1104 26682 38272 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38272 26682
rect 1104 26608 38272 26630
rect 6914 26528 6920 26580
rect 6972 26568 6978 26580
rect 7745 26571 7803 26577
rect 7745 26568 7757 26571
rect 6972 26540 7757 26568
rect 6972 26528 6978 26540
rect 7745 26537 7757 26540
rect 7791 26537 7803 26571
rect 7745 26531 7803 26537
rect 7944 26540 8340 26568
rect 7944 26500 7972 26540
rect 7392 26472 7972 26500
rect 8312 26500 8340 26540
rect 12250 26528 12256 26580
rect 12308 26568 12314 26580
rect 13446 26568 13452 26580
rect 12308 26540 13452 26568
rect 12308 26528 12314 26540
rect 13446 26528 13452 26540
rect 13504 26528 13510 26580
rect 13817 26571 13875 26577
rect 13817 26537 13829 26571
rect 13863 26568 13875 26571
rect 14274 26568 14280 26580
rect 13863 26540 14280 26568
rect 13863 26537 13875 26540
rect 13817 26531 13875 26537
rect 14274 26528 14280 26540
rect 14332 26528 14338 26580
rect 14461 26571 14519 26577
rect 14461 26537 14473 26571
rect 14507 26568 14519 26571
rect 14642 26568 14648 26580
rect 14507 26540 14648 26568
rect 14507 26537 14519 26540
rect 14461 26531 14519 26537
rect 14642 26528 14648 26540
rect 14700 26528 14706 26580
rect 17310 26568 17316 26580
rect 15028 26540 17316 26568
rect 11238 26500 11244 26512
rect 8312 26472 11244 26500
rect 7282 26432 7288 26444
rect 4540 26404 7288 26432
rect 4540 26373 4568 26404
rect 7282 26392 7288 26404
rect 7340 26392 7346 26444
rect 7392 26373 7420 26472
rect 11238 26460 11244 26472
rect 11296 26460 11302 26512
rect 14918 26500 14924 26512
rect 12406 26472 14924 26500
rect 7561 26435 7619 26441
rect 7561 26401 7573 26435
rect 7607 26432 7619 26435
rect 7834 26432 7840 26444
rect 7607 26404 7840 26432
rect 7607 26401 7619 26404
rect 7561 26395 7619 26401
rect 7834 26392 7840 26404
rect 7892 26392 7898 26444
rect 8110 26392 8116 26444
rect 8168 26432 8174 26444
rect 8665 26435 8723 26441
rect 8665 26432 8677 26435
rect 8168 26404 8677 26432
rect 8168 26392 8174 26404
rect 8665 26401 8677 26404
rect 8711 26432 8723 26435
rect 8754 26432 8760 26444
rect 8711 26404 8760 26432
rect 8711 26401 8723 26404
rect 8665 26395 8723 26401
rect 8754 26392 8760 26404
rect 8812 26392 8818 26444
rect 12406 26432 12434 26472
rect 14918 26460 14924 26472
rect 14976 26460 14982 26512
rect 8864 26404 12434 26432
rect 4525 26367 4583 26373
rect 4525 26333 4537 26367
rect 4571 26333 4583 26367
rect 4525 26327 4583 26333
rect 4617 26367 4675 26373
rect 4617 26333 4629 26367
rect 4663 26364 4675 26367
rect 4801 26367 4859 26373
rect 4801 26364 4813 26367
rect 4663 26336 4813 26364
rect 4663 26333 4675 26336
rect 4617 26327 4675 26333
rect 4801 26333 4813 26336
rect 4847 26333 4859 26367
rect 4801 26327 4859 26333
rect 7377 26367 7435 26373
rect 7377 26333 7389 26367
rect 7423 26333 7435 26367
rect 7377 26327 7435 26333
rect 7929 26367 7987 26373
rect 7929 26333 7941 26367
rect 7975 26333 7987 26367
rect 7929 26327 7987 26333
rect 5074 26256 5080 26308
rect 5132 26256 5138 26308
rect 6825 26299 6883 26305
rect 5460 26268 5566 26296
rect 3878 26188 3884 26240
rect 3936 26228 3942 26240
rect 5460 26228 5488 26268
rect 6825 26265 6837 26299
rect 6871 26296 6883 26299
rect 6871 26268 7328 26296
rect 6871 26265 6883 26268
rect 6825 26259 6883 26265
rect 5994 26228 6000 26240
rect 3936 26200 6000 26228
rect 3936 26188 3942 26200
rect 5994 26188 6000 26200
rect 6052 26188 6058 26240
rect 6914 26188 6920 26240
rect 6972 26188 6978 26240
rect 7300 26237 7328 26268
rect 7285 26231 7343 26237
rect 7285 26197 7297 26231
rect 7331 26228 7343 26231
rect 7834 26228 7840 26240
rect 7331 26200 7840 26228
rect 7331 26197 7343 26200
rect 7285 26191 7343 26197
rect 7834 26188 7840 26200
rect 7892 26188 7898 26240
rect 7944 26228 7972 26327
rect 8386 26324 8392 26376
rect 8444 26324 8450 26376
rect 8864 26364 8892 26404
rect 12894 26392 12900 26444
rect 12952 26432 12958 26444
rect 12952 26404 13584 26432
rect 12952 26392 12958 26404
rect 8588 26336 8892 26364
rect 9125 26367 9183 26373
rect 8478 26256 8484 26308
rect 8536 26256 8542 26308
rect 8021 26231 8079 26237
rect 8021 26228 8033 26231
rect 7944 26200 8033 26228
rect 8021 26197 8033 26200
rect 8067 26197 8079 26231
rect 8021 26191 8079 26197
rect 8110 26188 8116 26240
rect 8168 26228 8174 26240
rect 8588 26228 8616 26336
rect 9125 26333 9137 26367
rect 9171 26364 9183 26367
rect 9582 26364 9588 26376
rect 9171 26336 9588 26364
rect 9171 26333 9183 26336
rect 9125 26327 9183 26333
rect 9582 26324 9588 26336
rect 9640 26324 9646 26376
rect 11882 26324 11888 26376
rect 11940 26364 11946 26376
rect 12618 26364 12624 26376
rect 11940 26336 12624 26364
rect 11940 26324 11946 26336
rect 12618 26324 12624 26336
rect 12676 26324 12682 26376
rect 13556 26373 13584 26404
rect 14274 26392 14280 26444
rect 14332 26432 14338 26444
rect 14332 26404 14688 26432
rect 14332 26392 14338 26404
rect 13541 26367 13599 26373
rect 13541 26333 13553 26367
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 13630 26324 13636 26376
rect 13688 26324 13694 26376
rect 13909 26367 13967 26373
rect 13909 26333 13921 26367
rect 13955 26364 13967 26367
rect 13998 26364 14004 26376
rect 13955 26336 14004 26364
rect 13955 26333 13967 26336
rect 13909 26327 13967 26333
rect 13998 26324 14004 26336
rect 14056 26324 14062 26376
rect 14660 26373 14688 26404
rect 15028 26373 15056 26540
rect 17310 26528 17316 26540
rect 17368 26528 17374 26580
rect 17405 26571 17463 26577
rect 17405 26537 17417 26571
rect 17451 26568 17463 26571
rect 17678 26568 17684 26580
rect 17451 26540 17684 26568
rect 17451 26537 17463 26540
rect 17405 26531 17463 26537
rect 17678 26528 17684 26540
rect 17736 26528 17742 26580
rect 18598 26528 18604 26580
rect 18656 26568 18662 26580
rect 19150 26568 19156 26580
rect 18656 26540 19156 26568
rect 18656 26528 18662 26540
rect 19150 26528 19156 26540
rect 19208 26528 19214 26580
rect 25406 26568 25412 26580
rect 19306 26540 25412 26568
rect 15102 26460 15108 26512
rect 15160 26460 15166 26512
rect 15562 26460 15568 26512
rect 15620 26460 15626 26512
rect 17862 26500 17868 26512
rect 17420 26472 17868 26500
rect 15470 26432 15476 26444
rect 15212 26404 15476 26432
rect 14645 26367 14703 26373
rect 14645 26333 14657 26367
rect 14691 26333 14703 26367
rect 14645 26327 14703 26333
rect 15013 26367 15071 26373
rect 15013 26333 15025 26367
rect 15059 26333 15071 26367
rect 15013 26327 15071 26333
rect 13357 26299 13415 26305
rect 13357 26265 13369 26299
rect 13403 26296 13415 26299
rect 14550 26296 14556 26308
rect 13403 26268 14556 26296
rect 13403 26265 13415 26268
rect 13357 26259 13415 26265
rect 14550 26256 14556 26268
rect 14608 26256 14614 26308
rect 14737 26299 14795 26305
rect 14737 26265 14749 26299
rect 14783 26265 14795 26299
rect 14737 26259 14795 26265
rect 14829 26299 14887 26305
rect 14829 26265 14841 26299
rect 14875 26296 14887 26299
rect 15212 26296 15240 26404
rect 15470 26392 15476 26404
rect 15528 26392 15534 26444
rect 15286 26324 15292 26376
rect 15344 26324 15350 26376
rect 15381 26367 15439 26373
rect 15381 26333 15393 26367
rect 15427 26364 15439 26367
rect 15580 26364 15608 26460
rect 15672 26404 17172 26432
rect 15672 26373 15700 26404
rect 15427 26336 15608 26364
rect 15657 26367 15715 26373
rect 15427 26333 15439 26336
rect 15381 26327 15439 26333
rect 15657 26333 15669 26367
rect 15703 26333 15715 26367
rect 15657 26327 15715 26333
rect 15746 26324 15752 26376
rect 15804 26364 15810 26376
rect 16209 26367 16267 26373
rect 16209 26364 16221 26367
rect 15804 26336 16221 26364
rect 15804 26324 15810 26336
rect 16209 26333 16221 26336
rect 16255 26333 16267 26367
rect 16209 26327 16267 26333
rect 16853 26367 16911 26373
rect 16853 26333 16865 26367
rect 16899 26364 16911 26367
rect 16942 26364 16948 26376
rect 16899 26336 16948 26364
rect 16899 26333 16911 26336
rect 16853 26327 16911 26333
rect 16942 26324 16948 26336
rect 17000 26324 17006 26376
rect 14875 26268 15240 26296
rect 14875 26265 14887 26268
rect 14829 26259 14887 26265
rect 8168 26200 8616 26228
rect 8168 26188 8174 26200
rect 8662 26188 8668 26240
rect 8720 26228 8726 26240
rect 9033 26231 9091 26237
rect 9033 26228 9045 26231
rect 8720 26200 9045 26228
rect 8720 26188 8726 26200
rect 9033 26197 9045 26200
rect 9079 26197 9091 26231
rect 9033 26191 9091 26197
rect 12342 26188 12348 26240
rect 12400 26228 12406 26240
rect 14752 26228 14780 26259
rect 15470 26256 15476 26308
rect 15528 26256 15534 26308
rect 15764 26228 15792 26324
rect 15930 26256 15936 26308
rect 15988 26296 15994 26308
rect 17144 26305 17172 26404
rect 17267 26367 17325 26373
rect 17267 26333 17279 26367
rect 17313 26364 17325 26367
rect 17420 26364 17448 26472
rect 17862 26460 17868 26472
rect 17920 26460 17926 26512
rect 17954 26460 17960 26512
rect 18012 26500 18018 26512
rect 19306 26500 19334 26540
rect 18012 26472 19334 26500
rect 21361 26503 21419 26509
rect 18012 26460 18018 26472
rect 21361 26469 21373 26503
rect 21407 26500 21419 26503
rect 22646 26500 22652 26512
rect 21407 26472 22652 26500
rect 21407 26469 21419 26472
rect 21361 26463 21419 26469
rect 22646 26460 22652 26472
rect 22704 26460 22710 26512
rect 17770 26392 17776 26444
rect 17828 26432 17834 26444
rect 25332 26432 25360 26540
rect 25406 26528 25412 26540
rect 25464 26528 25470 26580
rect 25498 26528 25504 26580
rect 25556 26568 25562 26580
rect 27801 26571 27859 26577
rect 25556 26540 25820 26568
rect 25556 26528 25562 26540
rect 17828 26404 24624 26432
rect 25332 26404 25452 26432
rect 17828 26392 17834 26404
rect 17313 26336 17448 26364
rect 17313 26333 17325 26336
rect 17267 26327 17325 26333
rect 17494 26324 17500 26376
rect 17552 26364 17558 26376
rect 20806 26364 20812 26376
rect 17552 26336 20812 26364
rect 17552 26324 17558 26336
rect 20806 26324 20812 26336
rect 20864 26324 20870 26376
rect 20898 26324 20904 26376
rect 20956 26364 20962 26376
rect 21085 26367 21143 26373
rect 21085 26364 21097 26367
rect 20956 26336 21097 26364
rect 20956 26324 20962 26336
rect 21085 26333 21097 26336
rect 21131 26333 21143 26367
rect 21085 26327 21143 26333
rect 21177 26367 21235 26373
rect 21177 26333 21189 26367
rect 21223 26333 21235 26367
rect 21177 26327 21235 26333
rect 16025 26299 16083 26305
rect 16025 26296 16037 26299
rect 15988 26268 16037 26296
rect 15988 26256 15994 26268
rect 16025 26265 16037 26268
rect 16071 26265 16083 26299
rect 16025 26259 16083 26265
rect 16393 26299 16451 26305
rect 16393 26265 16405 26299
rect 16439 26296 16451 26299
rect 17037 26299 17095 26305
rect 17037 26296 17049 26299
rect 16439 26268 17049 26296
rect 16439 26265 16451 26268
rect 16393 26259 16451 26265
rect 17037 26265 17049 26268
rect 17083 26265 17095 26299
rect 17037 26259 17095 26265
rect 17129 26299 17187 26305
rect 17129 26265 17141 26299
rect 17175 26265 17187 26299
rect 17129 26259 17187 26265
rect 12400 26200 15792 26228
rect 17144 26228 17172 26259
rect 17678 26256 17684 26308
rect 17736 26296 17742 26308
rect 20162 26296 20168 26308
rect 17736 26268 20168 26296
rect 17736 26256 17742 26268
rect 20162 26256 20168 26268
rect 20220 26296 20226 26308
rect 20257 26299 20315 26305
rect 20257 26296 20269 26299
rect 20220 26268 20269 26296
rect 20220 26256 20226 26268
rect 20257 26265 20269 26268
rect 20303 26265 20315 26299
rect 20257 26259 20315 26265
rect 20438 26256 20444 26308
rect 20496 26256 20502 26308
rect 20625 26299 20683 26305
rect 20625 26265 20637 26299
rect 20671 26296 20683 26299
rect 20993 26299 21051 26305
rect 20993 26296 21005 26299
rect 20671 26268 21005 26296
rect 20671 26265 20683 26268
rect 20625 26259 20683 26265
rect 20993 26265 21005 26268
rect 21039 26265 21051 26299
rect 21192 26296 21220 26327
rect 22922 26324 22928 26376
rect 22980 26364 22986 26376
rect 23290 26364 23296 26376
rect 22980 26336 23296 26364
rect 22980 26324 22986 26336
rect 23290 26324 23296 26336
rect 23348 26364 23354 26376
rect 23569 26367 23627 26373
rect 23569 26364 23581 26367
rect 23348 26336 23581 26364
rect 23348 26324 23354 26336
rect 23569 26333 23581 26336
rect 23615 26333 23627 26367
rect 23569 26327 23627 26333
rect 23845 26367 23903 26373
rect 23845 26333 23857 26367
rect 23891 26364 23903 26367
rect 24486 26364 24492 26376
rect 23891 26336 24492 26364
rect 23891 26333 23903 26336
rect 23845 26327 23903 26333
rect 24486 26324 24492 26336
rect 24544 26324 24550 26376
rect 21542 26296 21548 26308
rect 21192 26268 21548 26296
rect 20993 26259 21051 26265
rect 21542 26256 21548 26268
rect 21600 26256 21606 26308
rect 24596 26296 24624 26404
rect 24670 26324 24676 26376
rect 24728 26364 24734 26376
rect 25314 26364 25320 26376
rect 24728 26336 25320 26364
rect 24728 26324 24734 26336
rect 25314 26324 25320 26336
rect 25372 26324 25378 26376
rect 25424 26373 25452 26404
rect 25409 26367 25467 26373
rect 25409 26333 25421 26367
rect 25455 26333 25467 26367
rect 25409 26327 25467 26333
rect 25590 26324 25596 26376
rect 25648 26324 25654 26376
rect 25792 26373 25820 26540
rect 25884 26540 26924 26568
rect 25777 26367 25835 26373
rect 25777 26333 25789 26367
rect 25823 26333 25835 26367
rect 25777 26327 25835 26333
rect 25685 26299 25743 26305
rect 25685 26296 25697 26299
rect 24596 26268 25697 26296
rect 25685 26265 25697 26268
rect 25731 26296 25743 26299
rect 25884 26296 25912 26540
rect 25961 26503 26019 26509
rect 25961 26469 25973 26503
rect 26007 26469 26019 26503
rect 25961 26463 26019 26469
rect 25976 26432 26004 26463
rect 26142 26460 26148 26512
rect 26200 26500 26206 26512
rect 26896 26500 26924 26540
rect 27801 26537 27813 26571
rect 27847 26568 27859 26571
rect 28166 26568 28172 26580
rect 27847 26540 28172 26568
rect 27847 26537 27859 26540
rect 27801 26531 27859 26537
rect 28166 26528 28172 26540
rect 28224 26528 28230 26580
rect 30006 26528 30012 26580
rect 30064 26568 30070 26580
rect 30285 26571 30343 26577
rect 30285 26568 30297 26571
rect 30064 26540 30297 26568
rect 30064 26528 30070 26540
rect 30285 26537 30297 26540
rect 30331 26537 30343 26571
rect 30285 26531 30343 26537
rect 33134 26528 33140 26580
rect 33192 26568 33198 26580
rect 33229 26571 33287 26577
rect 33229 26568 33241 26571
rect 33192 26540 33241 26568
rect 33192 26528 33198 26540
rect 33229 26537 33241 26540
rect 33275 26537 33287 26571
rect 33229 26531 33287 26537
rect 29270 26500 29276 26512
rect 26200 26472 26832 26500
rect 26896 26472 29276 26500
rect 26200 26460 26206 26472
rect 25976 26404 26556 26432
rect 26050 26324 26056 26376
rect 26108 26324 26114 26376
rect 26234 26324 26240 26376
rect 26292 26324 26298 26376
rect 26528 26373 26556 26404
rect 26694 26392 26700 26444
rect 26752 26392 26758 26444
rect 26804 26432 26832 26472
rect 29270 26460 29276 26472
rect 29328 26460 29334 26512
rect 34885 26503 34943 26509
rect 29656 26472 30144 26500
rect 28258 26432 28264 26444
rect 26804 26404 28264 26432
rect 28258 26392 28264 26404
rect 28316 26392 28322 26444
rect 28350 26392 28356 26444
rect 28408 26432 28414 26444
rect 29656 26441 29684 26472
rect 30116 26444 30144 26472
rect 34885 26469 34897 26503
rect 34931 26469 34943 26503
rect 34885 26463 34943 26469
rect 29641 26435 29699 26441
rect 29641 26432 29653 26435
rect 28408 26404 29653 26432
rect 28408 26392 28414 26404
rect 29641 26401 29653 26404
rect 29687 26401 29699 26435
rect 29641 26395 29699 26401
rect 30098 26392 30104 26444
rect 30156 26392 30162 26444
rect 30926 26432 30932 26444
rect 30392 26404 30932 26432
rect 26329 26367 26387 26373
rect 26329 26333 26341 26367
rect 26375 26333 26387 26367
rect 26329 26327 26387 26333
rect 26513 26367 26571 26373
rect 26513 26333 26525 26367
rect 26559 26333 26571 26367
rect 26513 26327 26571 26333
rect 26605 26367 26663 26373
rect 26605 26333 26617 26367
rect 26651 26364 26663 26367
rect 26712 26364 26740 26392
rect 28994 26364 29000 26376
rect 26651 26336 26740 26364
rect 26804 26336 29000 26364
rect 26651 26333 26663 26336
rect 26605 26327 26663 26333
rect 25731 26268 25912 26296
rect 26068 26296 26096 26324
rect 26344 26296 26372 26327
rect 26804 26296 26832 26336
rect 28994 26324 29000 26336
rect 29052 26364 29058 26376
rect 29825 26367 29883 26373
rect 29825 26364 29837 26367
rect 29052 26336 29837 26364
rect 29052 26324 29058 26336
rect 29825 26333 29837 26336
rect 29871 26333 29883 26367
rect 29825 26327 29883 26333
rect 30006 26324 30012 26376
rect 30064 26364 30070 26376
rect 30392 26364 30420 26404
rect 30926 26392 30932 26404
rect 30984 26392 30990 26444
rect 31297 26435 31355 26441
rect 31297 26401 31309 26435
rect 31343 26432 31355 26435
rect 31386 26432 31392 26444
rect 31343 26404 31392 26432
rect 31343 26401 31355 26404
rect 31297 26395 31355 26401
rect 31386 26392 31392 26404
rect 31444 26392 31450 26444
rect 32490 26392 32496 26444
rect 32548 26432 32554 26444
rect 33045 26435 33103 26441
rect 33045 26432 33057 26435
rect 32548 26404 33057 26432
rect 32548 26392 32554 26404
rect 33045 26401 33057 26404
rect 33091 26401 33103 26435
rect 33045 26395 33103 26401
rect 33870 26392 33876 26444
rect 33928 26392 33934 26444
rect 34900 26432 34928 26463
rect 35253 26435 35311 26441
rect 35253 26432 35265 26435
rect 34900 26404 35265 26432
rect 35253 26401 35265 26404
rect 35299 26401 35311 26435
rect 35253 26395 35311 26401
rect 30064 26336 30420 26364
rect 30064 26324 30070 26336
rect 30466 26324 30472 26376
rect 30524 26364 30530 26376
rect 30745 26367 30803 26373
rect 30745 26364 30757 26367
rect 30524 26336 30757 26364
rect 30524 26324 30530 26336
rect 30745 26333 30757 26336
rect 30791 26333 30803 26367
rect 30745 26327 30803 26333
rect 30837 26367 30895 26373
rect 30837 26333 30849 26367
rect 30883 26364 30895 26367
rect 31021 26367 31079 26373
rect 31021 26364 31033 26367
rect 30883 26336 31033 26364
rect 30883 26333 30895 26336
rect 30837 26327 30895 26333
rect 31021 26333 31033 26336
rect 31067 26333 31079 26367
rect 31021 26327 31079 26333
rect 32674 26324 32680 26376
rect 32732 26364 32738 26376
rect 33597 26367 33655 26373
rect 33597 26364 33609 26367
rect 32732 26336 33609 26364
rect 32732 26324 32738 26336
rect 33597 26333 33609 26336
rect 33643 26364 33655 26367
rect 33778 26364 33784 26376
rect 33643 26336 33784 26364
rect 33643 26333 33655 26336
rect 33597 26327 33655 26333
rect 33778 26324 33784 26336
rect 33836 26324 33842 26376
rect 34698 26324 34704 26376
rect 34756 26324 34762 26376
rect 34974 26324 34980 26376
rect 35032 26324 35038 26376
rect 28169 26299 28227 26305
rect 28169 26296 28181 26299
rect 26068 26268 26832 26296
rect 27356 26268 28181 26296
rect 25731 26265 25743 26268
rect 25685 26259 25743 26265
rect 27356 26240 27384 26268
rect 28169 26265 28181 26268
rect 28215 26265 28227 26299
rect 28169 26259 28227 26265
rect 29178 26256 29184 26308
rect 29236 26296 29242 26308
rect 29917 26299 29975 26305
rect 29917 26296 29929 26299
rect 29236 26268 29929 26296
rect 29236 26256 29242 26268
rect 29917 26265 29929 26268
rect 29963 26296 29975 26299
rect 31294 26296 31300 26308
rect 29963 26268 31300 26296
rect 29963 26265 29975 26268
rect 29917 26259 29975 26265
rect 31294 26256 31300 26268
rect 31352 26256 31358 26308
rect 31570 26256 31576 26308
rect 31628 26296 31634 26308
rect 31628 26268 31786 26296
rect 31628 26256 31634 26268
rect 32766 26256 32772 26308
rect 32824 26296 32830 26308
rect 33689 26299 33747 26305
rect 33689 26296 33701 26299
rect 32824 26268 33701 26296
rect 32824 26256 32830 26268
rect 33689 26265 33701 26268
rect 33735 26296 33747 26299
rect 34238 26296 34244 26308
rect 33735 26268 34244 26296
rect 33735 26265 33747 26268
rect 33689 26259 33747 26265
rect 34238 26256 34244 26268
rect 34296 26256 34302 26308
rect 35986 26256 35992 26308
rect 36044 26256 36050 26308
rect 36630 26256 36636 26308
rect 36688 26296 36694 26308
rect 37001 26299 37059 26305
rect 37001 26296 37013 26299
rect 36688 26268 37013 26296
rect 36688 26256 36694 26268
rect 37001 26265 37013 26268
rect 37047 26265 37059 26299
rect 37001 26259 37059 26265
rect 17310 26228 17316 26240
rect 17144 26200 17316 26228
rect 12400 26188 12406 26200
rect 17310 26188 17316 26200
rect 17368 26188 17374 26240
rect 20070 26188 20076 26240
rect 20128 26228 20134 26240
rect 22738 26228 22744 26240
rect 20128 26200 22744 26228
rect 20128 26188 20134 26200
rect 22738 26188 22744 26200
rect 22796 26188 22802 26240
rect 23382 26188 23388 26240
rect 23440 26188 23446 26240
rect 23750 26188 23756 26240
rect 23808 26188 23814 26240
rect 26050 26188 26056 26240
rect 26108 26188 26114 26240
rect 27338 26188 27344 26240
rect 27396 26188 27402 26240
rect 27798 26188 27804 26240
rect 27856 26228 27862 26240
rect 32674 26228 32680 26240
rect 27856 26200 32680 26228
rect 27856 26188 27862 26200
rect 32674 26188 32680 26200
rect 32732 26228 32738 26240
rect 33318 26228 33324 26240
rect 32732 26200 33324 26228
rect 32732 26188 32738 26200
rect 33318 26188 33324 26200
rect 33376 26188 33382 26240
rect 1104 26138 38272 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38272 26138
rect 1104 26064 38272 26086
rect 5074 25984 5080 26036
rect 5132 26024 5138 26036
rect 5445 26027 5503 26033
rect 5445 26024 5457 26027
rect 5132 25996 5457 26024
rect 5132 25984 5138 25996
rect 5445 25993 5457 25996
rect 5491 25993 5503 26027
rect 5445 25987 5503 25993
rect 6914 25984 6920 26036
rect 6972 25984 6978 26036
rect 16393 26027 16451 26033
rect 16393 25993 16405 26027
rect 16439 26024 16451 26027
rect 19242 26024 19248 26036
rect 16439 25996 19248 26024
rect 16439 25993 16451 25996
rect 16393 25987 16451 25993
rect 19242 25984 19248 25996
rect 19300 25984 19306 26036
rect 19794 26024 19800 26036
rect 19444 25996 19800 26024
rect 3878 25956 3884 25968
rect 2976 25928 3884 25956
rect 2976 25900 3004 25928
rect 3878 25916 3884 25928
rect 3936 25956 3942 25968
rect 3936 25928 4094 25956
rect 3936 25916 3942 25928
rect 1762 25848 1768 25900
rect 1820 25848 1826 25900
rect 2958 25848 2964 25900
rect 3016 25848 3022 25900
rect 3050 25848 3056 25900
rect 3108 25848 3114 25900
rect 5629 25891 5687 25897
rect 5629 25857 5641 25891
rect 5675 25888 5687 25891
rect 6932 25888 6960 25984
rect 16758 25916 16764 25968
rect 16816 25956 16822 25968
rect 17770 25956 17776 25968
rect 16816 25928 17776 25956
rect 16816 25916 16822 25928
rect 17770 25916 17776 25928
rect 17828 25916 17834 25968
rect 18414 25956 18420 25968
rect 17880 25928 18420 25956
rect 5675 25860 6960 25888
rect 5675 25857 5687 25860
rect 5629 25851 5687 25857
rect 10042 25848 10048 25900
rect 10100 25848 10106 25900
rect 13814 25848 13820 25900
rect 13872 25888 13878 25900
rect 16209 25891 16267 25897
rect 16209 25888 16221 25891
rect 13872 25860 16221 25888
rect 13872 25848 13878 25860
rect 16209 25857 16221 25860
rect 16255 25857 16267 25891
rect 17880 25888 17908 25928
rect 18414 25916 18420 25928
rect 18472 25956 18478 25968
rect 19061 25959 19119 25965
rect 18472 25928 18828 25956
rect 18472 25916 18478 25928
rect 16209 25851 16267 25857
rect 16500 25860 17908 25888
rect 1854 25780 1860 25832
rect 1912 25820 1918 25832
rect 3329 25823 3387 25829
rect 3329 25820 3341 25823
rect 1912 25792 3341 25820
rect 1912 25780 1918 25792
rect 3329 25789 3341 25792
rect 3375 25789 3387 25823
rect 3329 25783 3387 25789
rect 3602 25780 3608 25832
rect 3660 25780 3666 25832
rect 8662 25780 8668 25832
rect 8720 25780 8726 25832
rect 8938 25780 8944 25832
rect 8996 25780 9002 25832
rect 14642 25780 14648 25832
rect 14700 25820 14706 25832
rect 16500 25820 16528 25860
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18322 25888 18328 25900
rect 18012 25860 18328 25888
rect 18012 25848 18018 25860
rect 18322 25848 18328 25860
rect 18380 25888 18386 25900
rect 18800 25897 18828 25928
rect 19061 25925 19073 25959
rect 19107 25956 19119 25959
rect 19444 25956 19472 25996
rect 19794 25984 19800 25996
rect 19852 25984 19858 26036
rect 20806 25984 20812 26036
rect 20864 26024 20870 26036
rect 21174 26024 21180 26036
rect 20864 25996 21180 26024
rect 20864 25984 20870 25996
rect 21174 25984 21180 25996
rect 21232 25984 21238 26036
rect 22462 25984 22468 26036
rect 22520 25984 22526 26036
rect 23750 25984 23756 26036
rect 23808 26024 23814 26036
rect 23937 26027 23995 26033
rect 23937 26024 23949 26027
rect 23808 25996 23949 26024
rect 23808 25984 23814 25996
rect 23937 25993 23949 25996
rect 23983 25993 23995 26027
rect 23937 25987 23995 25993
rect 24762 25984 24768 26036
rect 24820 26024 24826 26036
rect 24820 25996 25084 26024
rect 24820 25984 24826 25996
rect 19107 25928 19472 25956
rect 19521 25959 19579 25965
rect 19107 25925 19119 25928
rect 19061 25919 19119 25925
rect 19521 25925 19533 25959
rect 19567 25956 19579 25959
rect 19886 25956 19892 25968
rect 19567 25928 19892 25956
rect 19567 25925 19579 25928
rect 19521 25919 19579 25925
rect 19886 25916 19892 25928
rect 19944 25956 19950 25968
rect 20254 25956 20260 25968
rect 19944 25928 20260 25956
rect 19944 25916 19950 25928
rect 20254 25916 20260 25928
rect 20312 25916 20318 25968
rect 20530 25916 20536 25968
rect 20588 25956 20594 25968
rect 20625 25959 20683 25965
rect 20625 25956 20637 25959
rect 20588 25928 20637 25956
rect 20588 25916 20594 25928
rect 20625 25925 20637 25928
rect 20671 25925 20683 25959
rect 22480 25956 22508 25984
rect 23014 25956 23020 25968
rect 22480 25928 23020 25956
rect 20625 25919 20683 25925
rect 23014 25916 23020 25928
rect 23072 25956 23078 25968
rect 25056 25956 25084 25996
rect 25130 25984 25136 26036
rect 25188 26024 25194 26036
rect 25225 26027 25283 26033
rect 25225 26024 25237 26027
rect 25188 25996 25237 26024
rect 25188 25984 25194 25996
rect 25225 25993 25237 25996
rect 25271 25993 25283 26027
rect 25225 25987 25283 25993
rect 25314 25984 25320 26036
rect 25372 26024 25378 26036
rect 25372 25996 26004 26024
rect 25372 25984 25378 25996
rect 23072 25928 23428 25956
rect 23072 25916 23078 25928
rect 18693 25891 18751 25897
rect 18693 25888 18705 25891
rect 18380 25860 18705 25888
rect 18380 25848 18386 25860
rect 18693 25857 18705 25860
rect 18739 25857 18751 25891
rect 18693 25851 18751 25857
rect 18785 25891 18843 25897
rect 18785 25857 18797 25891
rect 18831 25857 18843 25891
rect 18785 25851 18843 25857
rect 18877 25891 18935 25897
rect 18877 25857 18889 25891
rect 18923 25888 18935 25891
rect 18966 25888 18972 25900
rect 18923 25860 18972 25888
rect 18923 25857 18935 25860
rect 18877 25851 18935 25857
rect 14700 25792 16528 25820
rect 14700 25780 14706 25792
rect 16574 25780 16580 25832
rect 16632 25820 16638 25832
rect 18138 25820 18144 25832
rect 16632 25792 18144 25820
rect 16632 25780 16638 25792
rect 18138 25780 18144 25792
rect 18196 25780 18202 25832
rect 18414 25780 18420 25832
rect 18472 25820 18478 25832
rect 18892 25820 18920 25851
rect 18966 25848 18972 25860
rect 19024 25848 19030 25900
rect 19334 25897 19340 25900
rect 19312 25891 19340 25897
rect 19312 25857 19324 25891
rect 19312 25851 19340 25857
rect 19334 25848 19340 25851
rect 19392 25848 19398 25900
rect 19429 25891 19487 25897
rect 19429 25857 19441 25891
rect 19475 25857 19487 25891
rect 19429 25851 19487 25857
rect 19676 25891 19734 25897
rect 19676 25857 19688 25891
rect 19722 25888 19734 25891
rect 19722 25857 19748 25888
rect 19676 25851 19748 25857
rect 18472 25792 18920 25820
rect 19444 25820 19472 25851
rect 19720 25820 19748 25851
rect 19794 25848 19800 25900
rect 19852 25848 19858 25900
rect 20438 25848 20444 25900
rect 20496 25848 20502 25900
rect 20717 25891 20775 25897
rect 20717 25857 20729 25891
rect 20763 25857 20775 25891
rect 20717 25851 20775 25857
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25888 20867 25891
rect 20990 25888 20996 25900
rect 20855 25860 20996 25888
rect 20855 25857 20867 25860
rect 20809 25851 20867 25857
rect 20070 25820 20076 25832
rect 19444 25792 19656 25820
rect 19720 25792 20076 25820
rect 18472 25780 18478 25792
rect 15102 25712 15108 25764
rect 15160 25752 15166 25764
rect 18509 25755 18567 25761
rect 18509 25752 18521 25755
rect 15160 25724 18521 25752
rect 15160 25712 15166 25724
rect 18509 25721 18521 25724
rect 18555 25752 18567 25755
rect 19518 25752 19524 25764
rect 18555 25724 19524 25752
rect 18555 25721 18567 25724
rect 18509 25715 18567 25721
rect 19518 25712 19524 25724
rect 19576 25712 19582 25764
rect 934 25644 940 25696
rect 992 25684 998 25696
rect 1489 25687 1547 25693
rect 1489 25684 1501 25687
rect 992 25656 1501 25684
rect 992 25644 998 25656
rect 1489 25653 1501 25656
rect 1535 25653 1547 25687
rect 1489 25647 1547 25653
rect 2866 25644 2872 25696
rect 2924 25644 2930 25696
rect 5074 25644 5080 25696
rect 5132 25644 5138 25696
rect 9674 25644 9680 25696
rect 9732 25684 9738 25696
rect 10413 25687 10471 25693
rect 10413 25684 10425 25687
rect 9732 25656 10425 25684
rect 9732 25644 9738 25656
rect 10413 25653 10425 25656
rect 10459 25684 10471 25687
rect 13078 25684 13084 25696
rect 10459 25656 13084 25684
rect 10459 25653 10471 25656
rect 10413 25647 10471 25653
rect 13078 25644 13084 25656
rect 13136 25644 13142 25696
rect 18138 25644 18144 25696
rect 18196 25684 18202 25696
rect 19058 25684 19064 25696
rect 18196 25656 19064 25684
rect 18196 25644 18202 25656
rect 19058 25644 19064 25656
rect 19116 25644 19122 25696
rect 19150 25644 19156 25696
rect 19208 25644 19214 25696
rect 19334 25644 19340 25696
rect 19392 25684 19398 25696
rect 19628 25684 19656 25792
rect 20070 25780 20076 25792
rect 20128 25780 20134 25832
rect 19702 25712 19708 25764
rect 19760 25752 19766 25764
rect 20732 25752 20760 25851
rect 20990 25848 20996 25860
rect 21048 25848 21054 25900
rect 22186 25848 22192 25900
rect 22244 25888 22250 25900
rect 22465 25891 22523 25897
rect 22465 25888 22477 25891
rect 22244 25860 22477 25888
rect 22244 25848 22250 25860
rect 22465 25857 22477 25860
rect 22511 25857 22523 25891
rect 22465 25851 22523 25857
rect 22646 25848 22652 25900
rect 22704 25848 22710 25900
rect 22741 25891 22799 25897
rect 22741 25857 22753 25891
rect 22787 25857 22799 25891
rect 22741 25851 22799 25857
rect 21008 25820 21036 25848
rect 21008 25792 22692 25820
rect 19760 25724 21128 25752
rect 19760 25712 19766 25724
rect 21100 25696 21128 25724
rect 22066 25724 22416 25752
rect 20898 25684 20904 25696
rect 19392 25656 20904 25684
rect 19392 25644 19398 25656
rect 20898 25644 20904 25656
rect 20956 25644 20962 25696
rect 20990 25644 20996 25696
rect 21048 25644 21054 25696
rect 21082 25644 21088 25696
rect 21140 25644 21146 25696
rect 21266 25644 21272 25696
rect 21324 25684 21330 25696
rect 22066 25684 22094 25724
rect 22388 25696 22416 25724
rect 22554 25712 22560 25764
rect 22612 25712 22618 25764
rect 21324 25656 22094 25684
rect 21324 25644 21330 25656
rect 22278 25644 22284 25696
rect 22336 25644 22342 25696
rect 22370 25644 22376 25696
rect 22428 25644 22434 25696
rect 22664 25684 22692 25792
rect 22756 25752 22784 25851
rect 23106 25848 23112 25900
rect 23164 25848 23170 25900
rect 23400 25897 23428 25928
rect 23768 25928 24992 25956
rect 25056 25928 25912 25956
rect 23385 25891 23443 25897
rect 23385 25857 23397 25891
rect 23431 25857 23443 25891
rect 23385 25851 23443 25857
rect 22922 25780 22928 25832
rect 22980 25820 22986 25832
rect 22980 25792 23612 25820
rect 22980 25780 22986 25792
rect 23477 25755 23535 25761
rect 23477 25752 23489 25755
rect 22756 25724 23489 25752
rect 23477 25721 23489 25724
rect 23523 25721 23535 25755
rect 23477 25715 23535 25721
rect 23106 25684 23112 25696
rect 22664 25656 23112 25684
rect 23106 25644 23112 25656
rect 23164 25644 23170 25696
rect 23584 25684 23612 25792
rect 23658 25780 23664 25832
rect 23716 25820 23722 25832
rect 23768 25829 23796 25928
rect 23845 25891 23903 25897
rect 23845 25857 23857 25891
rect 23891 25888 23903 25891
rect 24302 25888 24308 25900
rect 23891 25860 24308 25888
rect 23891 25857 23903 25860
rect 23845 25851 23903 25857
rect 24302 25848 24308 25860
rect 24360 25848 24366 25900
rect 24581 25891 24639 25897
rect 24581 25857 24593 25891
rect 24627 25888 24639 25891
rect 24670 25888 24676 25900
rect 24627 25860 24676 25888
rect 24627 25857 24639 25860
rect 24581 25851 24639 25857
rect 24670 25848 24676 25860
rect 24728 25848 24734 25900
rect 24762 25848 24768 25900
rect 24820 25848 24826 25900
rect 24964 25897 24992 25928
rect 24857 25891 24915 25897
rect 24857 25857 24869 25891
rect 24903 25857 24915 25891
rect 24857 25851 24915 25857
rect 24949 25891 25007 25897
rect 24949 25857 24961 25891
rect 24995 25888 25007 25891
rect 25130 25888 25136 25900
rect 24995 25860 25136 25888
rect 24995 25857 25007 25860
rect 24949 25851 25007 25857
rect 23753 25823 23811 25829
rect 23753 25820 23765 25823
rect 23716 25792 23765 25820
rect 23716 25780 23722 25792
rect 23753 25789 23765 25792
rect 23799 25789 23811 25823
rect 23753 25783 23811 25789
rect 23934 25780 23940 25832
rect 23992 25820 23998 25832
rect 24210 25820 24216 25832
rect 23992 25792 24216 25820
rect 23992 25780 23998 25792
rect 24210 25780 24216 25792
rect 24268 25780 24274 25832
rect 24320 25820 24348 25848
rect 24872 25820 24900 25851
rect 25130 25848 25136 25860
rect 25188 25848 25194 25900
rect 25498 25888 25504 25900
rect 25240 25860 25504 25888
rect 25240 25820 25268 25860
rect 25498 25848 25504 25860
rect 25556 25848 25562 25900
rect 25884 25897 25912 25928
rect 25976 25897 26004 25996
rect 26050 25984 26056 26036
rect 26108 25984 26114 26036
rect 29638 25984 29644 26036
rect 29696 26024 29702 26036
rect 30098 26024 30104 26036
rect 29696 25996 30104 26024
rect 29696 25984 29702 25996
rect 30098 25984 30104 25996
rect 30156 25984 30162 26036
rect 31294 25984 31300 26036
rect 31352 26024 31358 26036
rect 31352 25996 31524 26024
rect 31352 25984 31358 25996
rect 25593 25891 25651 25897
rect 25593 25857 25605 25891
rect 25639 25857 25651 25891
rect 25593 25851 25651 25857
rect 25685 25891 25743 25897
rect 25685 25857 25697 25891
rect 25731 25888 25743 25891
rect 25869 25891 25927 25897
rect 25731 25860 25820 25888
rect 25731 25857 25743 25860
rect 25685 25851 25743 25857
rect 24320 25792 24900 25820
rect 24964 25792 25268 25820
rect 24964 25764 24992 25792
rect 25406 25780 25412 25832
rect 25464 25820 25470 25832
rect 25608 25820 25636 25851
rect 25464 25792 25636 25820
rect 25464 25780 25470 25792
rect 24946 25712 24952 25764
rect 25004 25712 25010 25764
rect 25590 25712 25596 25764
rect 25648 25752 25654 25764
rect 25792 25752 25820 25860
rect 25869 25857 25881 25891
rect 25915 25857 25927 25891
rect 25869 25851 25927 25857
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25857 26019 25891
rect 26068 25888 26096 25984
rect 31386 25956 31392 25968
rect 26344 25928 31392 25956
rect 26344 25900 26372 25928
rect 31386 25916 31392 25928
rect 31444 25916 31450 25968
rect 31496 25956 31524 25996
rect 31570 25984 31576 26036
rect 31628 25984 31634 26036
rect 31662 25984 31668 26036
rect 31720 26024 31726 26036
rect 32125 26027 32183 26033
rect 32125 26024 32137 26027
rect 31720 25996 32137 26024
rect 31720 25984 31726 25996
rect 32125 25993 32137 25996
rect 32171 25993 32183 26027
rect 32125 25987 32183 25993
rect 32490 25984 32496 26036
rect 32548 26024 32554 26036
rect 32585 26027 32643 26033
rect 32585 26024 32597 26027
rect 32548 25996 32597 26024
rect 32548 25984 32554 25996
rect 32585 25993 32597 25996
rect 32631 25993 32643 26027
rect 32585 25987 32643 25993
rect 34330 25984 34336 26036
rect 34388 25984 34394 26036
rect 34698 25984 34704 26036
rect 34756 26024 34762 26036
rect 34793 26027 34851 26033
rect 34793 26024 34805 26027
rect 34756 25996 34805 26024
rect 34756 25984 34762 25996
rect 34793 25993 34805 25996
rect 34839 25993 34851 26027
rect 34793 25987 34851 25993
rect 34974 25984 34980 26036
rect 35032 26024 35038 26036
rect 35253 26027 35311 26033
rect 35253 26024 35265 26027
rect 35032 25996 35265 26024
rect 35032 25984 35038 25996
rect 35253 25993 35265 25996
rect 35299 25993 35311 26027
rect 35253 25987 35311 25993
rect 31941 25959 31999 25965
rect 31496 25928 31892 25956
rect 26145 25891 26203 25897
rect 26145 25888 26157 25891
rect 26068 25860 26157 25888
rect 25961 25851 26019 25857
rect 26145 25857 26157 25860
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 26237 25891 26295 25897
rect 26237 25857 26249 25891
rect 26283 25857 26295 25891
rect 26237 25851 26295 25857
rect 25884 25820 25912 25851
rect 26050 25820 26056 25832
rect 25884 25792 26056 25820
rect 26050 25780 26056 25792
rect 26108 25780 26114 25832
rect 26252 25820 26280 25851
rect 26326 25848 26332 25900
rect 26384 25848 26390 25900
rect 27154 25848 27160 25900
rect 27212 25888 27218 25900
rect 31481 25891 31539 25897
rect 31481 25888 31493 25891
rect 27212 25860 31493 25888
rect 27212 25848 27218 25860
rect 31481 25857 31493 25860
rect 31527 25857 31539 25891
rect 31481 25851 31539 25857
rect 31754 25848 31760 25900
rect 31812 25848 31818 25900
rect 31864 25888 31892 25928
rect 31941 25925 31953 25959
rect 31987 25956 31999 25959
rect 34348 25956 34376 25984
rect 31987 25928 32996 25956
rect 34348 25928 35112 25956
rect 31987 25925 31999 25928
rect 31941 25919 31999 25925
rect 32493 25891 32551 25897
rect 32493 25888 32505 25891
rect 31864 25860 32505 25888
rect 32493 25857 32505 25860
rect 32539 25888 32551 25891
rect 32766 25888 32772 25900
rect 32539 25860 32772 25888
rect 32539 25857 32551 25860
rect 32493 25851 32551 25857
rect 32766 25848 32772 25860
rect 32824 25848 32830 25900
rect 32968 25897 32996 25928
rect 32953 25891 33011 25897
rect 32953 25857 32965 25891
rect 32999 25857 33011 25891
rect 32953 25851 33011 25857
rect 33137 25891 33195 25897
rect 33137 25857 33149 25891
rect 33183 25857 33195 25891
rect 33137 25851 33195 25857
rect 26252 25792 26372 25820
rect 26344 25764 26372 25792
rect 28626 25780 28632 25832
rect 28684 25820 28690 25832
rect 30650 25820 30656 25832
rect 28684 25792 30656 25820
rect 28684 25780 28690 25792
rect 30650 25780 30656 25792
rect 30708 25780 30714 25832
rect 32674 25780 32680 25832
rect 32732 25780 32738 25832
rect 25958 25752 25964 25764
rect 25648 25724 25964 25752
rect 25648 25712 25654 25724
rect 25958 25712 25964 25724
rect 26016 25712 26022 25764
rect 26326 25712 26332 25764
rect 26384 25712 26390 25764
rect 23661 25687 23719 25693
rect 23661 25684 23673 25687
rect 23584 25656 23673 25684
rect 23661 25653 23673 25656
rect 23707 25684 23719 25687
rect 24118 25684 24124 25696
rect 23707 25656 24124 25684
rect 23707 25653 23719 25656
rect 23661 25647 23719 25653
rect 24118 25644 24124 25656
rect 24176 25644 24182 25696
rect 25314 25644 25320 25696
rect 25372 25644 25378 25696
rect 26602 25644 26608 25696
rect 26660 25644 26666 25696
rect 27522 25644 27528 25696
rect 27580 25684 27586 25696
rect 30006 25684 30012 25696
rect 27580 25656 30012 25684
rect 27580 25644 27586 25656
rect 30006 25644 30012 25656
rect 30064 25644 30070 25696
rect 30282 25644 30288 25696
rect 30340 25684 30346 25696
rect 33152 25684 33180 25851
rect 33226 25848 33232 25900
rect 33284 25848 33290 25900
rect 33318 25848 33324 25900
rect 33376 25848 33382 25900
rect 35084 25897 35112 25928
rect 34425 25891 34483 25897
rect 34425 25857 34437 25891
rect 34471 25857 34483 25891
rect 34425 25851 34483 25857
rect 35069 25891 35127 25897
rect 35069 25857 35081 25891
rect 35115 25888 35127 25891
rect 35161 25891 35219 25897
rect 35161 25888 35173 25891
rect 35115 25860 35173 25888
rect 35115 25857 35127 25860
rect 35069 25851 35127 25857
rect 35161 25857 35173 25860
rect 35207 25857 35219 25891
rect 35161 25851 35219 25857
rect 33336 25752 33364 25848
rect 34146 25780 34152 25832
rect 34204 25780 34210 25832
rect 34238 25780 34244 25832
rect 34296 25820 34302 25832
rect 34333 25823 34391 25829
rect 34333 25820 34345 25823
rect 34296 25792 34345 25820
rect 34296 25780 34302 25792
rect 34333 25789 34345 25792
rect 34379 25789 34391 25823
rect 34333 25783 34391 25789
rect 34440 25820 34468 25851
rect 36630 25848 36636 25900
rect 36688 25848 36694 25900
rect 36648 25820 36676 25848
rect 34440 25792 36676 25820
rect 34440 25752 34468 25792
rect 33336 25724 34468 25752
rect 34698 25712 34704 25764
rect 34756 25752 34762 25764
rect 34977 25755 35035 25761
rect 34977 25752 34989 25755
rect 34756 25724 34989 25752
rect 34756 25712 34762 25724
rect 34977 25721 34989 25724
rect 35023 25721 35035 25755
rect 34977 25715 35035 25721
rect 30340 25656 33180 25684
rect 33597 25687 33655 25693
rect 30340 25644 30346 25656
rect 33597 25653 33609 25687
rect 33643 25684 33655 25687
rect 34790 25684 34796 25696
rect 33643 25656 34796 25684
rect 33643 25653 33655 25656
rect 33597 25647 33655 25653
rect 34790 25644 34796 25656
rect 34848 25644 34854 25696
rect 1104 25594 38272 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38272 25594
rect 1104 25520 38272 25542
rect 3602 25440 3608 25492
rect 3660 25480 3666 25492
rect 3881 25483 3939 25489
rect 3881 25480 3893 25483
rect 3660 25452 3893 25480
rect 3660 25440 3666 25452
rect 3881 25449 3893 25452
rect 3927 25449 3939 25483
rect 3881 25443 3939 25449
rect 8938 25440 8944 25492
rect 8996 25480 9002 25492
rect 9033 25483 9091 25489
rect 9033 25480 9045 25483
rect 8996 25452 9045 25480
rect 8996 25440 9002 25452
rect 9033 25449 9045 25452
rect 9079 25449 9091 25483
rect 9033 25443 9091 25449
rect 9674 25440 9680 25492
rect 9732 25440 9738 25492
rect 12176 25452 12940 25480
rect 2133 25347 2191 25353
rect 2133 25313 2145 25347
rect 2179 25344 2191 25347
rect 2866 25344 2872 25356
rect 2179 25316 2872 25344
rect 2179 25313 2191 25316
rect 2133 25307 2191 25313
rect 2866 25304 2872 25316
rect 2924 25304 2930 25356
rect 1394 25236 1400 25288
rect 1452 25276 1458 25288
rect 1854 25276 1860 25288
rect 1452 25248 1860 25276
rect 1452 25236 1458 25248
rect 1854 25236 1860 25248
rect 1912 25236 1918 25288
rect 4065 25279 4123 25285
rect 4065 25245 4077 25279
rect 4111 25276 4123 25279
rect 4338 25276 4344 25288
rect 4111 25248 4344 25276
rect 4111 25245 4123 25248
rect 4065 25239 4123 25245
rect 4338 25236 4344 25248
rect 4396 25236 4402 25288
rect 7558 25236 7564 25288
rect 7616 25236 7622 25288
rect 9692 25285 9720 25440
rect 11885 25415 11943 25421
rect 11885 25381 11897 25415
rect 11931 25412 11943 25415
rect 12176 25412 12204 25452
rect 11931 25384 12204 25412
rect 11931 25381 11943 25384
rect 11885 25375 11943 25381
rect 9858 25304 9864 25356
rect 9916 25304 9922 25356
rect 9217 25279 9275 25285
rect 9217 25245 9229 25279
rect 9263 25276 9275 25279
rect 9677 25279 9735 25285
rect 9263 25248 9352 25276
rect 9263 25245 9275 25248
rect 9217 25239 9275 25245
rect 2866 25168 2872 25220
rect 2924 25168 2930 25220
rect 7576 25208 7604 25236
rect 9030 25208 9036 25220
rect 7576 25180 9036 25208
rect 9030 25168 9036 25180
rect 9088 25168 9094 25220
rect 3605 25143 3663 25149
rect 3605 25109 3617 25143
rect 3651 25140 3663 25143
rect 4614 25140 4620 25152
rect 3651 25112 4620 25140
rect 3651 25109 3663 25112
rect 3605 25103 3663 25109
rect 4614 25100 4620 25112
rect 4672 25100 4678 25152
rect 7282 25100 7288 25152
rect 7340 25140 7346 25152
rect 9324 25149 9352 25248
rect 9677 25245 9689 25279
rect 9723 25245 9735 25279
rect 9677 25239 9735 25245
rect 10134 25236 10140 25288
rect 10192 25236 10198 25288
rect 12176 25276 12204 25384
rect 12805 25415 12863 25421
rect 12805 25381 12817 25415
rect 12851 25381 12863 25415
rect 12912 25412 12940 25452
rect 13078 25440 13084 25492
rect 13136 25480 13142 25492
rect 19242 25480 19248 25492
rect 13136 25452 19248 25480
rect 13136 25440 13142 25452
rect 19242 25440 19248 25452
rect 19300 25480 19306 25492
rect 20438 25480 20444 25492
rect 19300 25452 20444 25480
rect 19300 25440 19306 25452
rect 20438 25440 20444 25452
rect 20496 25440 20502 25492
rect 22462 25480 22468 25492
rect 20824 25452 22468 25480
rect 15102 25412 15108 25424
rect 12912 25384 15108 25412
rect 12805 25375 12863 25381
rect 12250 25304 12256 25356
rect 12308 25344 12314 25356
rect 12529 25347 12587 25353
rect 12529 25344 12541 25347
rect 12308 25316 12541 25344
rect 12308 25304 12314 25316
rect 12529 25313 12541 25316
rect 12575 25313 12587 25347
rect 12820 25344 12848 25375
rect 13170 25344 13176 25356
rect 12820 25316 13176 25344
rect 12529 25307 12587 25313
rect 13170 25304 13176 25316
rect 13228 25304 13234 25356
rect 12345 25279 12403 25285
rect 12345 25276 12357 25279
rect 12176 25248 12357 25276
rect 12345 25245 12357 25248
rect 12391 25245 12403 25279
rect 12345 25239 12403 25245
rect 12618 25236 12624 25288
rect 12676 25276 12682 25288
rect 12943 25279 13001 25285
rect 12943 25276 12955 25279
rect 12676 25248 12955 25276
rect 12676 25236 12682 25248
rect 12943 25245 12955 25248
rect 12989 25245 13001 25279
rect 12943 25239 13001 25245
rect 13078 25236 13084 25288
rect 13136 25236 13142 25288
rect 13316 25285 13344 25384
rect 15102 25372 15108 25384
rect 15160 25372 15166 25424
rect 15194 25372 15200 25424
rect 15252 25412 15258 25424
rect 16393 25415 16451 25421
rect 16393 25412 16405 25415
rect 15252 25384 16405 25412
rect 15252 25372 15258 25384
rect 16393 25381 16405 25384
rect 16439 25381 16451 25415
rect 16393 25375 16451 25381
rect 17126 25372 17132 25424
rect 17184 25412 17190 25424
rect 17184 25384 17356 25412
rect 17184 25372 17190 25384
rect 14826 25304 14832 25356
rect 14884 25304 14890 25356
rect 15672 25316 17264 25344
rect 15672 25288 15700 25316
rect 13301 25279 13359 25285
rect 13301 25245 13313 25279
rect 13347 25245 13359 25279
rect 13301 25239 13359 25245
rect 13446 25236 13452 25288
rect 13504 25236 13510 25288
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25245 14611 25279
rect 14553 25239 14611 25245
rect 10413 25211 10471 25217
rect 10413 25177 10425 25211
rect 10459 25208 10471 25211
rect 10502 25208 10508 25220
rect 10459 25180 10508 25208
rect 10459 25177 10471 25180
rect 10413 25171 10471 25177
rect 10502 25168 10508 25180
rect 10560 25168 10566 25220
rect 11054 25168 11060 25220
rect 11112 25168 11118 25220
rect 11790 25168 11796 25220
rect 11848 25208 11854 25220
rect 12437 25211 12495 25217
rect 12437 25208 12449 25211
rect 11848 25180 12449 25208
rect 11848 25168 11854 25180
rect 12437 25177 12449 25180
rect 12483 25177 12495 25211
rect 12437 25171 12495 25177
rect 12526 25168 12532 25220
rect 12584 25208 12590 25220
rect 13173 25211 13231 25217
rect 13173 25208 13185 25211
rect 12584 25180 13185 25208
rect 12584 25168 12590 25180
rect 13173 25177 13185 25180
rect 13219 25208 13231 25211
rect 14182 25208 14188 25220
rect 13219 25180 14188 25208
rect 13219 25177 13231 25180
rect 13173 25171 13231 25177
rect 14182 25168 14188 25180
rect 14240 25208 14246 25220
rect 14568 25208 14596 25239
rect 15654 25236 15660 25288
rect 15712 25236 15718 25288
rect 15933 25279 15991 25285
rect 15933 25245 15945 25279
rect 15979 25276 15991 25279
rect 16206 25276 16212 25288
rect 15979 25248 16212 25276
rect 15979 25245 15991 25248
rect 15933 25239 15991 25245
rect 16206 25236 16212 25248
rect 16264 25236 16270 25288
rect 16761 25279 16819 25285
rect 16668 25257 16726 25263
rect 16668 25223 16680 25257
rect 16714 25223 16726 25257
rect 16761 25245 16773 25279
rect 16807 25245 16819 25279
rect 16761 25239 16819 25245
rect 16853 25279 16911 25285
rect 16853 25245 16865 25279
rect 16899 25276 16911 25279
rect 16942 25276 16948 25288
rect 16899 25248 16948 25276
rect 16899 25245 16911 25248
rect 16853 25239 16911 25245
rect 16668 25217 16726 25223
rect 14240 25180 14596 25208
rect 14240 25168 14246 25180
rect 7469 25143 7527 25149
rect 7469 25140 7481 25143
rect 7340 25112 7481 25140
rect 7340 25100 7346 25112
rect 7469 25109 7481 25112
rect 7515 25109 7527 25143
rect 7469 25103 7527 25109
rect 9309 25143 9367 25149
rect 9309 25109 9321 25143
rect 9355 25109 9367 25143
rect 9309 25103 9367 25109
rect 9582 25100 9588 25152
rect 9640 25140 9646 25152
rect 9769 25143 9827 25149
rect 9769 25140 9781 25143
rect 9640 25112 9781 25140
rect 9640 25100 9646 25112
rect 9769 25109 9781 25112
rect 9815 25140 9827 25143
rect 11808 25140 11836 25168
rect 9815 25112 11836 25140
rect 9815 25109 9827 25112
rect 9769 25103 9827 25109
rect 11974 25100 11980 25152
rect 12032 25100 12038 25152
rect 12342 25100 12348 25152
rect 12400 25140 12406 25152
rect 12802 25140 12808 25152
rect 12400 25112 12808 25140
rect 12400 25100 12406 25112
rect 12802 25100 12808 25112
rect 12860 25100 12866 25152
rect 16117 25143 16175 25149
rect 16117 25109 16129 25143
rect 16163 25140 16175 25143
rect 16683 25140 16711 25217
rect 16776 25208 16804 25239
rect 16942 25236 16948 25248
rect 17000 25236 17006 25288
rect 17034 25236 17040 25288
rect 17092 25236 17098 25288
rect 17236 25285 17264 25316
rect 17221 25279 17279 25285
rect 17221 25245 17233 25279
rect 17267 25245 17279 25279
rect 17221 25239 17279 25245
rect 17328 25208 17356 25384
rect 17862 25372 17868 25424
rect 17920 25412 17926 25424
rect 20824 25412 20852 25452
rect 22462 25440 22468 25452
rect 22520 25440 22526 25492
rect 22554 25440 22560 25492
rect 22612 25480 22618 25492
rect 22833 25483 22891 25489
rect 22833 25480 22845 25483
rect 22612 25452 22845 25480
rect 22612 25440 22618 25452
rect 22833 25449 22845 25452
rect 22879 25449 22891 25483
rect 22833 25443 22891 25449
rect 23566 25440 23572 25492
rect 23624 25440 23630 25492
rect 24762 25440 24768 25492
rect 24820 25440 24826 25492
rect 26878 25480 26884 25492
rect 24872 25452 26884 25480
rect 17920 25384 20852 25412
rect 17920 25372 17926 25384
rect 17405 25347 17463 25353
rect 17405 25313 17417 25347
rect 17451 25344 17463 25347
rect 18138 25344 18144 25356
rect 17451 25316 18144 25344
rect 17451 25313 17463 25316
rect 17405 25307 17463 25313
rect 18138 25304 18144 25316
rect 18196 25304 18202 25356
rect 19076 25353 19104 25384
rect 20898 25372 20904 25424
rect 20956 25412 20962 25424
rect 20956 25384 21128 25412
rect 20956 25372 20962 25384
rect 19061 25347 19119 25353
rect 19061 25313 19073 25347
rect 19107 25344 19119 25347
rect 19107 25316 19141 25344
rect 19107 25313 19119 25316
rect 19061 25307 19119 25313
rect 20990 25304 20996 25356
rect 21048 25304 21054 25356
rect 18230 25236 18236 25288
rect 18288 25276 18294 25288
rect 18325 25279 18383 25285
rect 18325 25276 18337 25279
rect 18288 25248 18337 25276
rect 18288 25236 18294 25248
rect 18325 25245 18337 25248
rect 18371 25245 18383 25279
rect 18325 25239 18383 25245
rect 18506 25236 18512 25288
rect 18564 25236 18570 25288
rect 18601 25279 18659 25285
rect 18601 25245 18613 25279
rect 18647 25245 18659 25279
rect 18601 25239 18659 25245
rect 18616 25208 18644 25239
rect 20714 25236 20720 25288
rect 20772 25236 20778 25288
rect 20901 25279 20959 25285
rect 20901 25245 20913 25279
rect 20947 25245 20959 25279
rect 20901 25239 20959 25245
rect 20070 25208 20076 25220
rect 16776 25180 17172 25208
rect 17328 25180 20076 25208
rect 17144 25152 17172 25180
rect 20070 25168 20076 25180
rect 20128 25208 20134 25220
rect 20346 25208 20352 25220
rect 20128 25180 20352 25208
rect 20128 25168 20134 25180
rect 20346 25168 20352 25180
rect 20404 25168 20410 25220
rect 16758 25140 16764 25152
rect 16163 25112 16764 25140
rect 16163 25109 16175 25112
rect 16117 25103 16175 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 17126 25100 17132 25152
rect 17184 25100 17190 25152
rect 17862 25100 17868 25152
rect 17920 25140 17926 25152
rect 19886 25140 19892 25152
rect 17920 25112 19892 25140
rect 17920 25100 17926 25112
rect 19886 25100 19892 25112
rect 19944 25100 19950 25152
rect 20533 25143 20591 25149
rect 20533 25109 20545 25143
rect 20579 25140 20591 25143
rect 20622 25140 20628 25152
rect 20579 25112 20628 25140
rect 20579 25109 20591 25112
rect 20533 25103 20591 25109
rect 20622 25100 20628 25112
rect 20680 25100 20686 25152
rect 20916 25140 20944 25239
rect 21100 25208 21128 25384
rect 21266 25372 21272 25424
rect 21324 25372 21330 25424
rect 21284 25344 21312 25372
rect 21284 25316 21404 25344
rect 21174 25236 21180 25288
rect 21232 25285 21238 25288
rect 21376 25285 21404 25316
rect 21232 25279 21281 25285
rect 21232 25245 21235 25279
rect 21269 25245 21281 25279
rect 21232 25239 21281 25245
rect 21361 25279 21419 25285
rect 21361 25245 21373 25279
rect 21407 25245 21419 25279
rect 21361 25239 21419 25245
rect 21232 25236 21238 25239
rect 21450 25236 21456 25288
rect 21508 25236 21514 25288
rect 21581 25279 21639 25285
rect 21581 25245 21593 25279
rect 21627 25245 21639 25279
rect 21581 25239 21639 25245
rect 21596 25208 21624 25239
rect 21726 25236 21732 25288
rect 21784 25236 21790 25288
rect 21836 25248 22140 25276
rect 21100 25180 21624 25208
rect 21085 25143 21143 25149
rect 21085 25140 21097 25143
rect 20916 25112 21097 25140
rect 21085 25109 21097 25112
rect 21131 25109 21143 25143
rect 21085 25103 21143 25109
rect 21174 25100 21180 25152
rect 21232 25140 21238 25152
rect 21836 25140 21864 25248
rect 22002 25168 22008 25220
rect 22060 25168 22066 25220
rect 22112 25208 22140 25248
rect 22186 25236 22192 25288
rect 22244 25236 22250 25288
rect 22370 25285 22376 25288
rect 22337 25279 22376 25285
rect 22337 25245 22349 25279
rect 22337 25239 22376 25245
rect 22370 25236 22376 25239
rect 22428 25236 22434 25288
rect 22480 25276 22508 25440
rect 22646 25372 22652 25424
rect 22704 25412 22710 25424
rect 23584 25412 23612 25440
rect 22704 25384 23612 25412
rect 22704 25372 22710 25384
rect 24210 25372 24216 25424
rect 24268 25412 24274 25424
rect 24872 25412 24900 25452
rect 26878 25440 26884 25452
rect 26936 25480 26942 25492
rect 31846 25480 31852 25492
rect 26936 25452 31852 25480
rect 26936 25440 26942 25452
rect 31846 25440 31852 25452
rect 31904 25480 31910 25492
rect 33318 25480 33324 25492
rect 31904 25452 33324 25480
rect 31904 25440 31910 25452
rect 33318 25440 33324 25452
rect 33376 25440 33382 25492
rect 26234 25412 26240 25424
rect 24268 25384 24900 25412
rect 24964 25384 26240 25412
rect 24268 25372 24274 25384
rect 23106 25304 23112 25356
rect 23164 25304 23170 25356
rect 23474 25304 23480 25356
rect 23532 25304 23538 25356
rect 22654 25279 22712 25285
rect 22654 25276 22666 25279
rect 22480 25248 22666 25276
rect 22654 25245 22666 25248
rect 22700 25245 22712 25279
rect 22654 25239 22712 25245
rect 23017 25279 23075 25285
rect 23017 25245 23029 25279
rect 23063 25245 23075 25279
rect 23124 25276 23152 25304
rect 24964 25285 24992 25384
rect 26234 25372 26240 25384
rect 26292 25372 26298 25424
rect 26418 25372 26424 25424
rect 26476 25372 26482 25424
rect 27801 25415 27859 25421
rect 27801 25381 27813 25415
rect 27847 25381 27859 25415
rect 27801 25375 27859 25381
rect 26142 25344 26148 25356
rect 25056 25316 26148 25344
rect 25056 25285 25084 25316
rect 26142 25304 26148 25316
rect 26200 25304 26206 25356
rect 26436 25344 26464 25372
rect 27522 25344 27528 25356
rect 26436 25316 27528 25344
rect 24949 25279 25007 25285
rect 24949 25276 24961 25279
rect 23124 25248 24961 25276
rect 23017 25239 23075 25245
rect 24949 25245 24961 25248
rect 24995 25245 25007 25279
rect 24949 25239 25007 25245
rect 25041 25279 25099 25285
rect 25041 25245 25053 25279
rect 25087 25245 25099 25279
rect 25041 25239 25099 25245
rect 25225 25279 25283 25285
rect 25225 25245 25237 25279
rect 25271 25245 25283 25279
rect 25225 25239 25283 25245
rect 25317 25279 25375 25285
rect 25317 25245 25329 25279
rect 25363 25276 25375 25279
rect 25363 25248 25452 25276
rect 25363 25245 25375 25248
rect 25317 25239 25375 25245
rect 22462 25208 22468 25220
rect 22112 25180 22468 25208
rect 22462 25168 22468 25180
rect 22520 25168 22526 25220
rect 22557 25211 22615 25217
rect 22557 25177 22569 25211
rect 22603 25177 22615 25211
rect 23032 25208 23060 25239
rect 22557 25171 22615 25177
rect 22664 25180 23060 25208
rect 21232 25112 21864 25140
rect 22020 25140 22048 25168
rect 22572 25140 22600 25171
rect 22664 25152 22692 25180
rect 22020 25112 22600 25140
rect 21232 25100 21238 25112
rect 22646 25100 22652 25152
rect 22704 25100 22710 25152
rect 22738 25100 22744 25152
rect 22796 25140 22802 25152
rect 25056 25140 25084 25239
rect 25240 25208 25268 25239
rect 25240 25180 25360 25208
rect 25332 25152 25360 25180
rect 22796 25112 25084 25140
rect 22796 25100 22802 25112
rect 25314 25100 25320 25152
rect 25372 25100 25378 25152
rect 25424 25140 25452 25248
rect 26050 25236 26056 25288
rect 26108 25236 26114 25288
rect 26786 25236 26792 25288
rect 26844 25276 26850 25288
rect 27448 25285 27476 25316
rect 27522 25304 27528 25316
rect 27580 25304 27586 25356
rect 27816 25344 27844 25375
rect 27890 25372 27896 25424
rect 27948 25412 27954 25424
rect 28902 25412 28908 25424
rect 27948 25384 28908 25412
rect 27948 25372 27954 25384
rect 28902 25372 28908 25384
rect 28960 25412 28966 25424
rect 28960 25384 30420 25412
rect 28960 25372 28966 25384
rect 27816 25316 28764 25344
rect 27157 25279 27215 25285
rect 27157 25276 27169 25279
rect 26844 25248 27169 25276
rect 26844 25236 26850 25248
rect 27157 25245 27169 25248
rect 27203 25245 27215 25279
rect 27157 25239 27215 25245
rect 27250 25279 27308 25285
rect 27250 25245 27262 25279
rect 27296 25245 27308 25279
rect 27250 25239 27308 25245
rect 27433 25279 27491 25285
rect 27433 25245 27445 25279
rect 27479 25245 27491 25279
rect 27433 25239 27491 25245
rect 27622 25279 27680 25285
rect 27622 25245 27634 25279
rect 27668 25245 27680 25279
rect 27622 25239 27680 25245
rect 26068 25208 26096 25236
rect 27265 25208 27293 25239
rect 26068 25180 27293 25208
rect 27522 25168 27528 25220
rect 27580 25168 27586 25220
rect 26694 25140 26700 25152
rect 25424 25112 26700 25140
rect 26694 25100 26700 25112
rect 26752 25100 26758 25152
rect 27154 25100 27160 25152
rect 27212 25140 27218 25152
rect 27632 25140 27660 25239
rect 28258 25236 28264 25288
rect 28316 25236 28322 25288
rect 28445 25279 28503 25285
rect 28445 25245 28457 25279
rect 28491 25276 28503 25279
rect 28626 25276 28632 25288
rect 28491 25248 28632 25276
rect 28491 25245 28503 25248
rect 28445 25239 28503 25245
rect 28626 25236 28632 25248
rect 28684 25236 28690 25288
rect 28736 25285 28764 25316
rect 29086 25304 29092 25356
rect 29144 25344 29150 25356
rect 29144 25316 29224 25344
rect 29144 25304 29150 25316
rect 29196 25285 29224 25316
rect 30116 25316 30328 25344
rect 28721 25279 28779 25285
rect 28721 25245 28733 25279
rect 28767 25245 28779 25279
rect 28721 25239 28779 25245
rect 29181 25279 29239 25285
rect 29181 25245 29193 25279
rect 29227 25245 29239 25279
rect 29181 25239 29239 25245
rect 30009 25279 30067 25285
rect 30009 25245 30021 25279
rect 30055 25245 30067 25279
rect 30009 25239 30067 25245
rect 28276 25208 28304 25236
rect 28537 25211 28595 25217
rect 28537 25208 28549 25211
rect 28276 25180 28549 25208
rect 28537 25177 28549 25180
rect 28583 25177 28595 25211
rect 28537 25171 28595 25177
rect 28905 25211 28963 25217
rect 28905 25177 28917 25211
rect 28951 25208 28963 25211
rect 30024 25208 30052 25239
rect 30116 25220 30144 25316
rect 30300 25285 30328 25316
rect 30392 25285 30420 25384
rect 34698 25372 34704 25424
rect 34756 25372 34762 25424
rect 30193 25279 30251 25285
rect 30193 25245 30205 25279
rect 30239 25245 30251 25279
rect 30193 25239 30251 25245
rect 30285 25279 30343 25285
rect 30285 25245 30297 25279
rect 30331 25245 30343 25279
rect 30285 25239 30343 25245
rect 30377 25279 30435 25285
rect 30377 25245 30389 25279
rect 30423 25276 30435 25279
rect 30926 25276 30932 25288
rect 30423 25248 30932 25276
rect 30423 25245 30435 25248
rect 30377 25239 30435 25245
rect 28951 25180 30052 25208
rect 28951 25177 28963 25180
rect 28905 25171 28963 25177
rect 30098 25168 30104 25220
rect 30156 25168 30162 25220
rect 30208 25208 30236 25239
rect 30926 25236 30932 25248
rect 30984 25236 30990 25288
rect 34330 25236 34336 25288
rect 34388 25236 34394 25288
rect 34716 25285 34744 25372
rect 34701 25279 34759 25285
rect 34701 25245 34713 25279
rect 34747 25245 34759 25279
rect 34701 25239 34759 25245
rect 34977 25211 35035 25217
rect 34977 25208 34989 25211
rect 30208 25180 30328 25208
rect 30300 25152 30328 25180
rect 34532 25180 34989 25208
rect 27212 25112 27660 25140
rect 27212 25100 27218 25112
rect 29086 25100 29092 25152
rect 29144 25100 29150 25152
rect 30282 25100 30288 25152
rect 30340 25100 30346 25152
rect 30653 25143 30711 25149
rect 30653 25109 30665 25143
rect 30699 25140 30711 25143
rect 31294 25140 31300 25152
rect 30699 25112 31300 25140
rect 30699 25109 30711 25112
rect 30653 25103 30711 25109
rect 31294 25100 31300 25112
rect 31352 25100 31358 25152
rect 34532 25149 34560 25180
rect 34977 25177 34989 25180
rect 35023 25177 35035 25211
rect 34977 25171 35035 25177
rect 35986 25168 35992 25220
rect 36044 25168 36050 25220
rect 36722 25168 36728 25220
rect 36780 25168 36786 25220
rect 34517 25143 34575 25149
rect 34517 25109 34529 25143
rect 34563 25109 34575 25143
rect 34517 25103 34575 25109
rect 1104 25050 38272 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38272 25050
rect 1104 24976 38272 24998
rect 4338 24896 4344 24948
rect 4396 24896 4402 24948
rect 4709 24939 4767 24945
rect 4709 24905 4721 24939
rect 4755 24936 4767 24939
rect 5074 24936 5080 24948
rect 4755 24908 5080 24936
rect 4755 24905 4767 24908
rect 4709 24899 4767 24905
rect 5074 24896 5080 24908
rect 5132 24936 5138 24948
rect 5810 24936 5816 24948
rect 5132 24908 5816 24936
rect 5132 24896 5138 24908
rect 5810 24896 5816 24908
rect 5868 24896 5874 24948
rect 9214 24896 9220 24948
rect 9272 24896 9278 24948
rect 9582 24896 9588 24948
rect 9640 24896 9646 24948
rect 10134 24896 10140 24948
rect 10192 24936 10198 24948
rect 10321 24939 10379 24945
rect 10321 24936 10333 24939
rect 10192 24908 10333 24936
rect 10192 24896 10198 24908
rect 10321 24905 10333 24908
rect 10367 24905 10379 24939
rect 10321 24899 10379 24905
rect 10502 24896 10508 24948
rect 10560 24936 10566 24948
rect 10597 24939 10655 24945
rect 10597 24936 10609 24939
rect 10560 24908 10609 24936
rect 10560 24896 10566 24908
rect 10597 24905 10609 24908
rect 10643 24905 10655 24939
rect 10597 24899 10655 24905
rect 11974 24896 11980 24948
rect 12032 24896 12038 24948
rect 12713 24939 12771 24945
rect 12713 24905 12725 24939
rect 12759 24936 12771 24939
rect 12759 24908 12848 24936
rect 12759 24905 12771 24908
rect 12713 24899 12771 24905
rect 5994 24828 6000 24880
rect 6052 24868 6058 24880
rect 6052 24840 8050 24868
rect 6052 24828 6058 24840
rect 2806 24772 2912 24800
rect 2884 24744 2912 24772
rect 5902 24760 5908 24812
rect 5960 24760 5966 24812
rect 10410 24760 10416 24812
rect 10468 24760 10474 24812
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24800 10839 24803
rect 11992 24800 12020 24896
rect 12342 24828 12348 24880
rect 12400 24828 12406 24880
rect 12820 24877 12848 24908
rect 14182 24896 14188 24948
rect 14240 24936 14246 24948
rect 14277 24939 14335 24945
rect 14277 24936 14289 24939
rect 14240 24908 14289 24936
rect 14240 24896 14246 24908
rect 14277 24905 14289 24908
rect 14323 24905 14335 24939
rect 15194 24936 15200 24948
rect 14277 24899 14335 24905
rect 14384 24908 15200 24936
rect 12805 24871 12863 24877
rect 12805 24837 12817 24871
rect 12851 24837 12863 24871
rect 12805 24831 12863 24837
rect 12989 24871 13047 24877
rect 12989 24837 13001 24871
rect 13035 24868 13047 24871
rect 13170 24868 13176 24880
rect 13035 24840 13176 24868
rect 13035 24837 13047 24840
rect 12989 24831 13047 24837
rect 13170 24828 13176 24840
rect 13228 24828 13234 24880
rect 14384 24868 14412 24908
rect 15194 24896 15200 24908
rect 15252 24896 15258 24948
rect 16942 24896 16948 24948
rect 17000 24936 17006 24948
rect 17000 24908 17448 24936
rect 17000 24896 17006 24908
rect 14200 24840 14412 24868
rect 10827 24772 12020 24800
rect 12161 24803 12219 24809
rect 10827 24769 10839 24772
rect 10781 24763 10839 24769
rect 12161 24769 12173 24803
rect 12207 24800 12219 24803
rect 12250 24800 12256 24812
rect 12207 24772 12256 24800
rect 12207 24769 12219 24772
rect 12161 24763 12219 24769
rect 12250 24760 12256 24772
rect 12308 24760 12314 24812
rect 12437 24803 12495 24809
rect 12437 24769 12449 24803
rect 12483 24769 12495 24803
rect 12437 24763 12495 24769
rect 12529 24803 12587 24809
rect 12529 24769 12541 24803
rect 12575 24800 12587 24803
rect 13538 24800 13544 24812
rect 12575 24772 12756 24800
rect 12575 24769 12587 24772
rect 12529 24763 12587 24769
rect 1394 24692 1400 24744
rect 1452 24692 1458 24744
rect 1670 24692 1676 24744
rect 1728 24692 1734 24744
rect 2866 24692 2872 24744
rect 2924 24692 2930 24744
rect 4798 24692 4804 24744
rect 4856 24692 4862 24744
rect 4985 24735 5043 24741
rect 4985 24701 4997 24735
rect 5031 24701 5043 24735
rect 4985 24695 5043 24701
rect 3142 24556 3148 24608
rect 3200 24556 3206 24608
rect 3970 24556 3976 24608
rect 4028 24596 4034 24608
rect 5000 24596 5028 24695
rect 7282 24692 7288 24744
rect 7340 24692 7346 24744
rect 7561 24735 7619 24741
rect 7561 24701 7573 24735
rect 7607 24732 7619 24735
rect 7926 24732 7932 24744
rect 7607 24704 7932 24732
rect 7607 24701 7619 24704
rect 7561 24695 7619 24701
rect 7926 24692 7932 24704
rect 7984 24692 7990 24744
rect 9677 24735 9735 24741
rect 9677 24701 9689 24735
rect 9723 24732 9735 24735
rect 9723 24704 9757 24732
rect 9723 24701 9735 24704
rect 9677 24695 9735 24701
rect 9033 24667 9091 24673
rect 9033 24633 9045 24667
rect 9079 24664 9091 24667
rect 9692 24664 9720 24695
rect 9858 24692 9864 24744
rect 9916 24692 9922 24744
rect 12452 24732 12480 24763
rect 12728 24732 12756 24772
rect 13004 24772 13544 24800
rect 13004 24732 13032 24772
rect 13538 24760 13544 24772
rect 13596 24800 13602 24812
rect 14200 24800 14228 24840
rect 14550 24828 14556 24880
rect 14608 24868 14614 24880
rect 15746 24868 15752 24880
rect 14608 24840 15752 24868
rect 14608 24828 14614 24840
rect 15746 24828 15752 24840
rect 15804 24828 15810 24880
rect 16209 24871 16267 24877
rect 16209 24837 16221 24871
rect 16255 24868 16267 24871
rect 16298 24868 16304 24880
rect 16255 24840 16304 24868
rect 16255 24837 16267 24840
rect 16209 24831 16267 24837
rect 16298 24828 16304 24840
rect 16356 24828 16362 24880
rect 16758 24868 16764 24880
rect 16684 24840 16764 24868
rect 13596 24772 14228 24800
rect 14369 24803 14427 24809
rect 13596 24760 13602 24772
rect 14369 24769 14381 24803
rect 14415 24800 14427 24803
rect 14829 24803 14887 24809
rect 14415 24772 14596 24800
rect 14415 24769 14427 24772
rect 14369 24763 14427 24769
rect 14568 24744 14596 24772
rect 14829 24769 14841 24803
rect 14875 24769 14887 24803
rect 14829 24763 14887 24769
rect 9968 24704 12664 24732
rect 12728 24704 13032 24732
rect 9968 24664 9996 24704
rect 9079 24636 9996 24664
rect 9079 24633 9091 24636
rect 9033 24627 9091 24633
rect 4028 24568 5028 24596
rect 4028 24556 4034 24568
rect 5626 24556 5632 24608
rect 5684 24596 5690 24608
rect 5721 24599 5779 24605
rect 5721 24596 5733 24599
rect 5684 24568 5733 24596
rect 5684 24556 5690 24568
rect 5721 24565 5733 24568
rect 5767 24565 5779 24599
rect 5721 24559 5779 24565
rect 7098 24556 7104 24608
rect 7156 24596 7162 24608
rect 12526 24596 12532 24608
rect 7156 24568 12532 24596
rect 7156 24556 7162 24568
rect 12526 24556 12532 24568
rect 12584 24556 12590 24608
rect 12636 24596 12664 24704
rect 14550 24692 14556 24744
rect 14608 24692 14614 24744
rect 14734 24692 14740 24744
rect 14792 24732 14798 24744
rect 14844 24732 14872 24763
rect 15378 24760 15384 24812
rect 15436 24760 15442 24812
rect 16684 24809 16712 24840
rect 16758 24828 16764 24840
rect 16816 24868 16822 24880
rect 17420 24868 17448 24908
rect 17586 24896 17592 24948
rect 17644 24936 17650 24948
rect 18509 24939 18567 24945
rect 17644 24908 18460 24936
rect 17644 24896 17650 24908
rect 17678 24868 17684 24880
rect 16816 24840 17355 24868
rect 17420 24840 17684 24868
rect 16816 24828 16822 24840
rect 16669 24803 16727 24809
rect 16669 24769 16681 24803
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 16853 24803 16911 24809
rect 16853 24769 16865 24803
rect 16899 24800 16911 24803
rect 17126 24800 17132 24812
rect 16899 24772 17132 24800
rect 16899 24769 16911 24772
rect 16853 24763 16911 24769
rect 17126 24760 17132 24772
rect 17184 24760 17190 24812
rect 17221 24803 17279 24809
rect 17221 24769 17233 24803
rect 17267 24769 17279 24803
rect 17327 24800 17355 24840
rect 17678 24828 17684 24840
rect 17736 24828 17742 24880
rect 18230 24828 18236 24880
rect 18288 24868 18294 24880
rect 18325 24871 18383 24877
rect 18325 24868 18337 24871
rect 18288 24840 18337 24868
rect 18288 24828 18294 24840
rect 18325 24837 18337 24840
rect 18371 24837 18383 24871
rect 18432 24868 18460 24908
rect 18509 24905 18521 24939
rect 18555 24936 18567 24939
rect 18598 24936 18604 24948
rect 18555 24908 18604 24936
rect 18555 24905 18567 24908
rect 18509 24899 18567 24905
rect 18598 24896 18604 24908
rect 18656 24896 18662 24948
rect 18693 24939 18751 24945
rect 18693 24905 18705 24939
rect 18739 24905 18751 24939
rect 18693 24899 18751 24905
rect 18708 24868 18736 24899
rect 18874 24896 18880 24948
rect 18932 24936 18938 24948
rect 21269 24939 21327 24945
rect 21269 24936 21281 24939
rect 18932 24908 21281 24936
rect 18932 24896 18938 24908
rect 21269 24905 21281 24908
rect 21315 24936 21327 24939
rect 22922 24936 22928 24948
rect 21315 24908 22928 24936
rect 21315 24905 21327 24908
rect 21269 24899 21327 24905
rect 22922 24896 22928 24908
rect 22980 24896 22986 24948
rect 23014 24896 23020 24948
rect 23072 24936 23078 24948
rect 23385 24939 23443 24945
rect 23385 24936 23397 24939
rect 23072 24908 23397 24936
rect 23072 24896 23078 24908
rect 23385 24905 23397 24908
rect 23431 24905 23443 24939
rect 27433 24939 27491 24945
rect 27433 24936 27445 24939
rect 23385 24899 23443 24905
rect 25424 24908 27445 24936
rect 25424 24880 25452 24908
rect 27433 24905 27445 24908
rect 27479 24936 27491 24939
rect 27522 24936 27528 24948
rect 27479 24908 27528 24936
rect 27479 24905 27491 24908
rect 27433 24899 27491 24905
rect 27522 24896 27528 24908
rect 27580 24896 27586 24948
rect 29086 24896 29092 24948
rect 29144 24896 29150 24948
rect 30098 24896 30104 24948
rect 30156 24936 30162 24948
rect 33226 24936 33232 24948
rect 30156 24908 33232 24936
rect 30156 24896 30162 24908
rect 20990 24868 20996 24880
rect 18432 24840 20996 24868
rect 18325 24831 18383 24837
rect 20990 24828 20996 24840
rect 21048 24828 21054 24880
rect 21082 24828 21088 24880
rect 21140 24828 21146 24880
rect 21453 24871 21511 24877
rect 21453 24868 21465 24871
rect 21192 24840 21465 24868
rect 19794 24800 19800 24812
rect 17327 24772 19800 24800
rect 17221 24763 17279 24769
rect 14792 24704 14872 24732
rect 14792 24692 14798 24704
rect 14918 24692 14924 24744
rect 14976 24732 14982 24744
rect 15013 24735 15071 24741
rect 15013 24732 15025 24735
rect 14976 24704 15025 24732
rect 14976 24692 14982 24704
rect 15013 24701 15025 24704
rect 15059 24701 15071 24735
rect 15013 24695 15071 24701
rect 12912 24636 15240 24664
rect 12912 24596 12940 24636
rect 12636 24568 12940 24596
rect 13170 24556 13176 24608
rect 13228 24556 13234 24608
rect 14090 24556 14096 24608
rect 14148 24596 14154 24608
rect 15102 24596 15108 24608
rect 14148 24568 15108 24596
rect 14148 24556 14154 24568
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 15212 24596 15240 24636
rect 16850 24624 16856 24676
rect 16908 24664 16914 24676
rect 17236 24664 17264 24763
rect 19794 24760 19800 24772
rect 19852 24760 19858 24812
rect 20070 24760 20076 24812
rect 20128 24800 20134 24812
rect 21192 24800 21220 24840
rect 21453 24837 21465 24840
rect 21499 24837 21511 24871
rect 21453 24831 21511 24837
rect 22002 24828 22008 24880
rect 22060 24868 22066 24880
rect 25406 24868 25412 24880
rect 22060 24840 25412 24868
rect 22060 24828 22066 24840
rect 25406 24828 25412 24840
rect 25464 24828 25470 24880
rect 26418 24828 26424 24880
rect 26476 24868 26482 24880
rect 27338 24868 27344 24880
rect 26476 24840 27344 24868
rect 26476 24828 26482 24840
rect 27338 24828 27344 24840
rect 27396 24828 27402 24880
rect 29104 24868 29132 24896
rect 28920 24840 29132 24868
rect 20128 24772 21220 24800
rect 21361 24803 21419 24809
rect 20128 24760 20134 24772
rect 21361 24769 21373 24803
rect 21407 24800 21419 24803
rect 21542 24800 21548 24812
rect 21407 24772 21548 24800
rect 21407 24769 21419 24772
rect 21361 24763 21419 24769
rect 21542 24760 21548 24772
rect 21600 24760 21606 24812
rect 21726 24760 21732 24812
rect 21784 24800 21790 24812
rect 22646 24800 22652 24812
rect 21784 24772 22652 24800
rect 21784 24760 21790 24772
rect 22646 24760 22652 24772
rect 22704 24760 22710 24812
rect 23474 24760 23480 24812
rect 23532 24760 23538 24812
rect 23566 24760 23572 24812
rect 23624 24760 23630 24812
rect 24029 24803 24087 24809
rect 24029 24769 24041 24803
rect 24075 24800 24087 24803
rect 25130 24800 25136 24812
rect 24075 24772 25136 24800
rect 24075 24769 24087 24772
rect 24029 24763 24087 24769
rect 25130 24760 25136 24772
rect 25188 24760 25194 24812
rect 25866 24760 25872 24812
rect 25924 24760 25930 24812
rect 26145 24803 26203 24809
rect 26145 24769 26157 24803
rect 26191 24800 26203 24803
rect 28629 24803 28687 24809
rect 26191 24772 27016 24800
rect 26191 24769 26203 24772
rect 26145 24763 26203 24769
rect 17313 24735 17371 24741
rect 17313 24701 17325 24735
rect 17359 24732 17371 24735
rect 17678 24732 17684 24744
rect 17359 24704 17684 24732
rect 17359 24701 17371 24704
rect 17313 24695 17371 24701
rect 17678 24692 17684 24704
rect 17736 24692 17742 24744
rect 17862 24692 17868 24744
rect 17920 24692 17926 24744
rect 20438 24732 20444 24744
rect 17972 24704 20444 24732
rect 17972 24676 18000 24704
rect 20438 24692 20444 24704
rect 20496 24692 20502 24744
rect 21637 24735 21695 24741
rect 21637 24701 21649 24735
rect 21683 24732 21695 24735
rect 22186 24732 22192 24744
rect 21683 24704 22192 24732
rect 21683 24701 21695 24704
rect 21637 24695 21695 24701
rect 22186 24692 22192 24704
rect 22244 24692 22250 24744
rect 23584 24732 23612 24760
rect 23842 24732 23848 24744
rect 23584 24704 23848 24732
rect 23842 24692 23848 24704
rect 23900 24732 23906 24744
rect 24121 24735 24179 24741
rect 24121 24732 24133 24735
rect 23900 24704 24133 24732
rect 23900 24692 23906 24704
rect 24121 24701 24133 24704
rect 24167 24701 24179 24735
rect 24121 24695 24179 24701
rect 25406 24692 25412 24744
rect 25464 24732 25470 24744
rect 25777 24735 25835 24741
rect 25777 24732 25789 24735
rect 25464 24704 25789 24732
rect 25464 24692 25470 24704
rect 25777 24701 25789 24704
rect 25823 24701 25835 24735
rect 25777 24695 25835 24701
rect 17402 24664 17408 24676
rect 16908 24636 17408 24664
rect 16908 24624 16914 24636
rect 17402 24624 17408 24636
rect 17460 24664 17466 24676
rect 17954 24664 17960 24676
rect 17460 24636 17960 24664
rect 17460 24624 17466 24636
rect 17954 24624 17960 24636
rect 18012 24624 18018 24676
rect 19334 24664 19340 24676
rect 18432 24636 19340 24664
rect 18432 24596 18460 24636
rect 19334 24624 19340 24636
rect 19392 24624 19398 24676
rect 24210 24624 24216 24676
rect 24268 24664 24274 24676
rect 26988 24673 27016 24772
rect 28629 24769 28641 24803
rect 28675 24800 28687 24803
rect 28810 24800 28816 24812
rect 28675 24772 28816 24800
rect 28675 24769 28687 24772
rect 28629 24763 28687 24769
rect 28810 24760 28816 24772
rect 28868 24760 28874 24812
rect 28920 24809 28948 24840
rect 29638 24828 29644 24880
rect 29696 24828 29702 24880
rect 30926 24828 30932 24880
rect 30984 24828 30990 24880
rect 28905 24803 28963 24809
rect 28905 24769 28917 24803
rect 28951 24769 28963 24803
rect 28905 24763 28963 24769
rect 31110 24760 31116 24812
rect 31168 24760 31174 24812
rect 31588 24809 31616 24908
rect 33226 24896 33232 24908
rect 33284 24896 33290 24948
rect 33318 24896 33324 24948
rect 33376 24896 33382 24948
rect 34241 24939 34299 24945
rect 34241 24905 34253 24939
rect 34287 24936 34299 24939
rect 34330 24936 34336 24948
rect 34287 24908 34336 24936
rect 34287 24905 34299 24908
rect 34241 24899 34299 24905
rect 34330 24896 34336 24908
rect 34388 24896 34394 24948
rect 31846 24828 31852 24880
rect 31904 24828 31910 24880
rect 33336 24868 33364 24896
rect 34609 24871 34667 24877
rect 34609 24868 34621 24871
rect 33336 24840 34621 24868
rect 34609 24837 34621 24840
rect 34655 24868 34667 24871
rect 36722 24868 36728 24880
rect 34655 24840 36728 24868
rect 34655 24837 34667 24840
rect 34609 24831 34667 24837
rect 36722 24828 36728 24840
rect 36780 24828 36786 24880
rect 31297 24803 31355 24809
rect 31297 24769 31309 24803
rect 31343 24769 31355 24803
rect 31297 24763 31355 24769
rect 31573 24803 31631 24809
rect 31573 24769 31585 24803
rect 31619 24769 31631 24803
rect 31864 24800 31892 24828
rect 33045 24813 33103 24819
rect 31941 24803 31999 24809
rect 31941 24800 31953 24803
rect 31864 24772 31953 24800
rect 31573 24763 31631 24769
rect 31941 24769 31953 24772
rect 31987 24769 31999 24803
rect 33045 24800 33057 24813
rect 31941 24763 31999 24769
rect 32968 24779 33057 24800
rect 33091 24779 33103 24813
rect 32968 24773 33103 24779
rect 33229 24803 33287 24809
rect 32968 24772 33088 24773
rect 27525 24735 27583 24741
rect 27525 24701 27537 24735
rect 27571 24732 27583 24735
rect 27798 24732 27804 24744
rect 27571 24704 27804 24732
rect 27571 24701 27583 24704
rect 27525 24695 27583 24701
rect 26973 24667 27031 24673
rect 24268 24636 26096 24664
rect 24268 24624 24274 24636
rect 15212 24568 18460 24596
rect 18506 24556 18512 24608
rect 18564 24556 18570 24608
rect 19518 24556 19524 24608
rect 19576 24596 19582 24608
rect 21266 24596 21272 24608
rect 19576 24568 21272 24596
rect 19576 24556 19582 24568
rect 21266 24556 21272 24568
rect 21324 24556 21330 24608
rect 21358 24556 21364 24608
rect 21416 24596 21422 24608
rect 25498 24596 25504 24608
rect 21416 24568 25504 24596
rect 21416 24556 21422 24568
rect 25498 24556 25504 24568
rect 25556 24556 25562 24608
rect 25958 24556 25964 24608
rect 26016 24556 26022 24608
rect 26068 24596 26096 24636
rect 26973 24633 26985 24667
rect 27019 24633 27031 24667
rect 26973 24627 27031 24633
rect 27540 24596 27568 24695
rect 27798 24692 27804 24704
rect 27856 24692 27862 24744
rect 29181 24735 29239 24741
rect 29181 24732 29193 24735
rect 28828 24704 29193 24732
rect 28828 24673 28856 24704
rect 29181 24701 29193 24704
rect 29227 24701 29239 24735
rect 29181 24695 29239 24701
rect 29730 24692 29736 24744
rect 29788 24732 29794 24744
rect 31312 24732 31340 24763
rect 29788 24704 31340 24732
rect 32968 24732 32996 24772
rect 33229 24769 33241 24803
rect 33275 24800 33287 24803
rect 33505 24803 33563 24809
rect 33505 24800 33517 24803
rect 33275 24772 33517 24800
rect 33275 24769 33287 24772
rect 33229 24763 33287 24769
rect 33505 24769 33517 24772
rect 33551 24800 33563 24803
rect 33778 24800 33784 24812
rect 33551 24772 33784 24800
rect 33551 24769 33563 24772
rect 33505 24763 33563 24769
rect 33042 24732 33048 24744
rect 32968 24704 33048 24732
rect 29788 24692 29794 24704
rect 30300 24676 30328 24704
rect 33042 24692 33048 24704
rect 33100 24692 33106 24744
rect 33134 24692 33140 24744
rect 33192 24732 33198 24744
rect 33244 24732 33272 24763
rect 33778 24760 33784 24772
rect 33836 24760 33842 24812
rect 33192 24704 33272 24732
rect 33192 24692 33198 24704
rect 33318 24692 33324 24744
rect 33376 24732 33382 24744
rect 33413 24735 33471 24741
rect 33413 24732 33425 24735
rect 33376 24704 33425 24732
rect 33376 24692 33382 24704
rect 33413 24701 33425 24704
rect 33459 24701 33471 24735
rect 33413 24695 33471 24701
rect 34701 24735 34759 24741
rect 34701 24701 34713 24735
rect 34747 24701 34759 24735
rect 34701 24695 34759 24701
rect 34793 24735 34851 24741
rect 34793 24701 34805 24735
rect 34839 24701 34851 24735
rect 34793 24695 34851 24701
rect 28813 24667 28871 24673
rect 28813 24633 28825 24667
rect 28859 24633 28871 24667
rect 28813 24627 28871 24633
rect 30282 24624 30288 24676
rect 30340 24624 30346 24676
rect 34716 24664 34744 24695
rect 31128 24636 31754 24664
rect 26068 24568 27568 24596
rect 28994 24556 29000 24608
rect 29052 24596 29058 24608
rect 30190 24596 30196 24608
rect 29052 24568 30196 24596
rect 29052 24556 29058 24568
rect 30190 24556 30196 24568
rect 30248 24596 30254 24608
rect 31128 24596 31156 24636
rect 30248 24568 31156 24596
rect 30248 24556 30254 24568
rect 31202 24556 31208 24608
rect 31260 24556 31266 24608
rect 31726 24596 31754 24636
rect 33060 24636 34744 24664
rect 33060 24596 33088 24636
rect 31726 24568 33088 24596
rect 33137 24599 33195 24605
rect 33137 24565 33149 24599
rect 33183 24596 33195 24599
rect 33318 24596 33324 24608
rect 33183 24568 33324 24596
rect 33183 24565 33195 24568
rect 33137 24559 33195 24565
rect 33318 24556 33324 24568
rect 33376 24556 33382 24608
rect 33410 24556 33416 24608
rect 33468 24596 33474 24608
rect 34146 24596 34152 24608
rect 33468 24568 34152 24596
rect 33468 24556 33474 24568
rect 34146 24556 34152 24568
rect 34204 24596 34210 24608
rect 34808 24596 34836 24695
rect 34204 24568 34836 24596
rect 34204 24556 34210 24568
rect 1104 24506 38272 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38272 24506
rect 1104 24432 38272 24454
rect 1670 24352 1676 24404
rect 1728 24392 1734 24404
rect 1765 24395 1823 24401
rect 1765 24392 1777 24395
rect 1728 24364 1777 24392
rect 1728 24352 1734 24364
rect 1765 24361 1777 24364
rect 1811 24361 1823 24395
rect 1765 24355 1823 24361
rect 3050 24352 3056 24404
rect 3108 24392 3114 24404
rect 3789 24395 3847 24401
rect 3789 24392 3801 24395
rect 3108 24364 3801 24392
rect 3108 24352 3114 24364
rect 3789 24361 3801 24364
rect 3835 24361 3847 24395
rect 3789 24355 3847 24361
rect 4062 24352 4068 24404
rect 4120 24392 4126 24404
rect 7834 24392 7840 24404
rect 4120 24364 7840 24392
rect 4120 24352 4126 24364
rect 7834 24352 7840 24364
rect 7892 24352 7898 24404
rect 7926 24352 7932 24404
rect 7984 24352 7990 24404
rect 9214 24352 9220 24404
rect 9272 24352 9278 24404
rect 13725 24395 13783 24401
rect 13725 24361 13737 24395
rect 13771 24361 13783 24395
rect 13725 24355 13783 24361
rect 13909 24395 13967 24401
rect 13909 24361 13921 24395
rect 13955 24392 13967 24395
rect 15378 24392 15384 24404
rect 13955 24364 15384 24392
rect 13955 24361 13967 24364
rect 13909 24355 13967 24361
rect 1394 24284 1400 24336
rect 1452 24324 1458 24336
rect 1452 24296 5304 24324
rect 1452 24284 1458 24296
rect 2961 24259 3019 24265
rect 2961 24225 2973 24259
rect 3007 24256 3019 24259
rect 3234 24256 3240 24268
rect 3007 24228 3240 24256
rect 3007 24225 3019 24228
rect 2961 24219 3019 24225
rect 3234 24216 3240 24228
rect 3292 24256 3298 24268
rect 3970 24256 3976 24268
rect 3292 24228 3976 24256
rect 3292 24216 3298 24228
rect 3970 24216 3976 24228
rect 4028 24256 4034 24268
rect 5276 24265 5304 24296
rect 4341 24259 4399 24265
rect 4341 24256 4353 24259
rect 4028 24228 4353 24256
rect 4028 24216 4034 24228
rect 4341 24225 4353 24228
rect 4387 24225 4399 24259
rect 4341 24219 4399 24225
rect 5261 24259 5319 24265
rect 5261 24225 5273 24259
rect 5307 24225 5319 24259
rect 5261 24219 5319 24225
rect 5537 24259 5595 24265
rect 5537 24225 5549 24259
rect 5583 24256 5595 24259
rect 5626 24256 5632 24268
rect 5583 24228 5632 24256
rect 5583 24225 5595 24228
rect 5537 24219 5595 24225
rect 5626 24216 5632 24228
rect 5684 24216 5690 24268
rect 9232 24256 9260 24352
rect 13740 24324 13768 24355
rect 15378 24352 15384 24364
rect 15436 24352 15442 24404
rect 15838 24352 15844 24404
rect 15896 24392 15902 24404
rect 15896 24364 17080 24392
rect 15896 24352 15902 24364
rect 14734 24324 14740 24336
rect 13740 24296 14740 24324
rect 14734 24284 14740 24296
rect 14792 24284 14798 24336
rect 15194 24284 15200 24336
rect 15252 24284 15258 24336
rect 15562 24284 15568 24336
rect 15620 24324 15626 24336
rect 16853 24327 16911 24333
rect 16853 24324 16865 24327
rect 15620 24296 16865 24324
rect 15620 24284 15626 24296
rect 16853 24293 16865 24296
rect 16899 24293 16911 24327
rect 16853 24287 16911 24293
rect 8128 24228 9260 24256
rect 1949 24191 2007 24197
rect 1949 24157 1961 24191
rect 1995 24188 2007 24191
rect 4157 24191 4215 24197
rect 1995 24160 2360 24188
rect 1995 24157 2007 24160
rect 1949 24151 2007 24157
rect 2332 24061 2360 24160
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 4614 24188 4620 24200
rect 4203 24160 4620 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4614 24148 4620 24160
rect 4672 24148 4678 24200
rect 8128 24197 8156 24228
rect 12710 24216 12716 24268
rect 12768 24216 12774 24268
rect 12989 24259 13047 24265
rect 12989 24225 13001 24259
rect 13035 24256 13047 24259
rect 13722 24256 13728 24268
rect 13035 24228 13728 24256
rect 13035 24225 13047 24228
rect 12989 24219 13047 24225
rect 13722 24216 13728 24228
rect 13780 24216 13786 24268
rect 13832 24228 14596 24256
rect 8113 24191 8171 24197
rect 8113 24157 8125 24191
rect 8159 24157 8171 24191
rect 8113 24151 8171 24157
rect 9122 24148 9128 24200
rect 9180 24148 9186 24200
rect 12728 24188 12756 24216
rect 12805 24191 12863 24197
rect 12805 24188 12817 24191
rect 12728 24160 12817 24188
rect 12805 24157 12817 24160
rect 12851 24157 12863 24191
rect 12805 24151 12863 24157
rect 2685 24123 2743 24129
rect 2685 24089 2697 24123
rect 2731 24120 2743 24123
rect 3142 24120 3148 24132
rect 2731 24092 3148 24120
rect 2731 24089 2743 24092
rect 2685 24083 2743 24089
rect 3142 24080 3148 24092
rect 3200 24080 3206 24132
rect 5994 24080 6000 24132
rect 6052 24080 6058 24132
rect 13541 24123 13599 24129
rect 13541 24089 13553 24123
rect 13587 24120 13599 24123
rect 13832 24120 13860 24228
rect 14277 24191 14335 24197
rect 14277 24188 14289 24191
rect 13587 24092 13860 24120
rect 13924 24160 14289 24188
rect 13587 24089 13599 24092
rect 13541 24083 13599 24089
rect 13924 24064 13952 24160
rect 14277 24157 14289 24160
rect 14323 24157 14335 24191
rect 14277 24151 14335 24157
rect 14568 24132 14596 24228
rect 14752 24197 14780 24284
rect 15286 24216 15292 24268
rect 15344 24256 15350 24268
rect 16393 24259 16451 24265
rect 16393 24256 16405 24259
rect 15344 24228 16405 24256
rect 15344 24216 15350 24228
rect 16393 24225 16405 24228
rect 16439 24225 16451 24259
rect 16393 24219 16451 24225
rect 16758 24216 16764 24268
rect 16816 24216 16822 24268
rect 17052 24256 17080 24364
rect 18322 24352 18328 24404
rect 18380 24392 18386 24404
rect 18601 24395 18659 24401
rect 18601 24392 18613 24395
rect 18380 24364 18613 24392
rect 18380 24352 18386 24364
rect 18601 24361 18613 24364
rect 18647 24361 18659 24395
rect 18601 24355 18659 24361
rect 18785 24395 18843 24401
rect 18785 24361 18797 24395
rect 18831 24392 18843 24395
rect 19150 24392 19156 24404
rect 18831 24364 19156 24392
rect 18831 24361 18843 24364
rect 18785 24355 18843 24361
rect 19150 24352 19156 24364
rect 19208 24352 19214 24404
rect 23658 24392 23664 24404
rect 19306 24364 23664 24392
rect 17126 24284 17132 24336
rect 17184 24324 17190 24336
rect 17310 24324 17316 24336
rect 17184 24296 17316 24324
rect 17184 24284 17190 24296
rect 17310 24284 17316 24296
rect 17368 24284 17374 24336
rect 17954 24324 17960 24336
rect 17512 24296 17960 24324
rect 17512 24256 17540 24296
rect 17954 24284 17960 24296
rect 18012 24284 18018 24336
rect 18141 24327 18199 24333
rect 18141 24293 18153 24327
rect 18187 24324 18199 24327
rect 18690 24324 18696 24336
rect 18187 24296 18696 24324
rect 18187 24293 18199 24296
rect 18141 24287 18199 24293
rect 18690 24284 18696 24296
rect 18748 24284 18754 24336
rect 19306 24324 19334 24364
rect 23658 24352 23664 24364
rect 23716 24352 23722 24404
rect 25406 24352 25412 24404
rect 25464 24352 25470 24404
rect 25498 24352 25504 24404
rect 25556 24392 25562 24404
rect 27341 24395 27399 24401
rect 25556 24364 27292 24392
rect 25556 24352 25562 24364
rect 18800 24296 19334 24324
rect 19889 24327 19947 24333
rect 17052 24228 17540 24256
rect 14737 24191 14795 24197
rect 14737 24157 14749 24191
rect 14783 24188 14795 24191
rect 14918 24188 14924 24200
rect 14783 24160 14924 24188
rect 14783 24157 14795 24160
rect 14737 24151 14795 24157
rect 14918 24148 14924 24160
rect 14976 24148 14982 24200
rect 15102 24148 15108 24200
rect 15160 24188 15166 24200
rect 15197 24191 15255 24197
rect 15197 24188 15209 24191
rect 15160 24160 15209 24188
rect 15160 24148 15166 24160
rect 15197 24157 15209 24160
rect 15243 24157 15255 24191
rect 15197 24151 15255 24157
rect 15749 24191 15807 24197
rect 15749 24157 15761 24191
rect 15795 24157 15807 24191
rect 15749 24151 15807 24157
rect 14550 24080 14556 24132
rect 14608 24120 14614 24132
rect 15010 24120 15016 24132
rect 14608 24092 15016 24120
rect 14608 24080 14614 24092
rect 15010 24080 15016 24092
rect 15068 24120 15074 24132
rect 15764 24120 15792 24151
rect 15838 24148 15844 24200
rect 15896 24188 15902 24200
rect 15933 24191 15991 24197
rect 15933 24188 15945 24191
rect 15896 24160 15945 24188
rect 15896 24148 15902 24160
rect 15933 24157 15945 24160
rect 15979 24157 15991 24191
rect 15933 24151 15991 24157
rect 16022 24148 16028 24200
rect 16080 24148 16086 24200
rect 16151 24191 16209 24197
rect 16151 24157 16163 24191
rect 16197 24188 16209 24191
rect 16776 24188 16804 24216
rect 17327 24197 17355 24228
rect 17095 24191 17153 24197
rect 17095 24188 17107 24191
rect 16197 24160 17107 24188
rect 16197 24157 16209 24160
rect 16151 24151 16209 24157
rect 17095 24157 17107 24160
rect 17141 24157 17153 24191
rect 17095 24151 17153 24157
rect 17221 24191 17279 24197
rect 17221 24157 17233 24191
rect 17267 24157 17279 24191
rect 17221 24151 17279 24157
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24157 17371 24191
rect 17313 24151 17371 24157
rect 16942 24120 16948 24132
rect 15068 24092 16948 24120
rect 15068 24080 15074 24092
rect 16942 24080 16948 24092
rect 17000 24080 17006 24132
rect 17236 24120 17264 24151
rect 17494 24148 17500 24200
rect 17552 24148 17558 24200
rect 17862 24148 17868 24200
rect 17920 24148 17926 24200
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24188 18199 24191
rect 18230 24188 18236 24200
rect 18187 24160 18236 24188
rect 18187 24157 18199 24160
rect 18141 24151 18199 24157
rect 18230 24148 18236 24160
rect 18288 24148 18294 24200
rect 18690 24148 18696 24200
rect 18748 24148 18754 24200
rect 17402 24120 17408 24132
rect 17236 24092 17408 24120
rect 17402 24080 17408 24092
rect 17460 24080 17466 24132
rect 18800 24120 18828 24296
rect 18892 24256 18920 24296
rect 19889 24293 19901 24327
rect 19935 24324 19947 24327
rect 20346 24324 20352 24336
rect 19935 24296 20352 24324
rect 19935 24293 19947 24296
rect 19889 24287 19947 24293
rect 20346 24284 20352 24296
rect 20404 24324 20410 24336
rect 20717 24327 20775 24333
rect 20717 24324 20729 24327
rect 20404 24296 20729 24324
rect 20404 24284 20410 24296
rect 20717 24293 20729 24296
rect 20763 24293 20775 24327
rect 20717 24287 20775 24293
rect 22094 24284 22100 24336
rect 22152 24284 22158 24336
rect 23566 24324 23572 24336
rect 23308 24296 23572 24324
rect 18892 24228 18966 24256
rect 18938 24197 18966 24228
rect 19150 24216 19156 24268
rect 19208 24256 19214 24268
rect 19208 24228 19748 24256
rect 19208 24216 19214 24228
rect 18923 24191 18981 24197
rect 18923 24157 18935 24191
rect 18969 24157 18981 24191
rect 18923 24151 18981 24157
rect 19058 24148 19064 24200
rect 19116 24148 19122 24200
rect 19426 24148 19432 24200
rect 19484 24188 19490 24200
rect 19720 24197 19748 24228
rect 19794 24216 19800 24268
rect 19852 24256 19858 24268
rect 22002 24256 22008 24268
rect 19852 24228 20024 24256
rect 19852 24216 19858 24228
rect 19996 24200 20024 24228
rect 20364 24228 22008 24256
rect 19521 24191 19579 24197
rect 19521 24188 19533 24191
rect 19484 24160 19533 24188
rect 19484 24148 19490 24160
rect 19521 24157 19533 24160
rect 19567 24157 19579 24191
rect 19521 24151 19579 24157
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24157 19763 24191
rect 19705 24151 19763 24157
rect 19978 24148 19984 24200
rect 20036 24188 20042 24200
rect 20364 24197 20392 24228
rect 22002 24216 22008 24228
rect 22060 24216 22066 24268
rect 22646 24216 22652 24268
rect 22704 24256 22710 24268
rect 23308 24265 23336 24296
rect 23566 24284 23572 24296
rect 23624 24324 23630 24336
rect 24670 24324 24676 24336
rect 23624 24296 24676 24324
rect 23624 24284 23630 24296
rect 24670 24284 24676 24296
rect 24728 24284 24734 24336
rect 25424 24324 25452 24352
rect 25424 24296 25636 24324
rect 25608 24265 25636 24296
rect 26970 24284 26976 24336
rect 27028 24284 27034 24336
rect 27264 24324 27292 24364
rect 27341 24361 27353 24395
rect 27387 24392 27399 24395
rect 27522 24392 27528 24404
rect 27387 24364 27528 24392
rect 27387 24361 27399 24364
rect 27341 24355 27399 24361
rect 27522 24352 27528 24364
rect 27580 24352 27586 24404
rect 31202 24352 31208 24404
rect 31260 24352 31266 24404
rect 31757 24395 31815 24401
rect 31757 24361 31769 24395
rect 31803 24361 31815 24395
rect 31757 24355 31815 24361
rect 32785 24364 34468 24392
rect 30098 24324 30104 24336
rect 27264 24296 30104 24324
rect 23293 24259 23351 24265
rect 23293 24256 23305 24259
rect 22704 24228 23305 24256
rect 22704 24216 22710 24228
rect 23293 24225 23305 24228
rect 23339 24225 23351 24259
rect 25593 24259 25651 24265
rect 23293 24219 23351 24225
rect 23492 24228 24808 24256
rect 23492 24200 23520 24228
rect 20349 24191 20407 24197
rect 20036 24160 20300 24188
rect 20036 24148 20042 24160
rect 17880 24092 18828 24120
rect 2317 24055 2375 24061
rect 2317 24021 2329 24055
rect 2363 24021 2375 24055
rect 2317 24015 2375 24021
rect 2774 24012 2780 24064
rect 2832 24012 2838 24064
rect 4249 24055 4307 24061
rect 4249 24021 4261 24055
rect 4295 24052 4307 24055
rect 4614 24052 4620 24064
rect 4295 24024 4620 24052
rect 4295 24021 4307 24024
rect 4249 24015 4307 24021
rect 4614 24012 4620 24024
rect 4672 24012 4678 24064
rect 6914 24012 6920 24064
rect 6972 24052 6978 24064
rect 7009 24055 7067 24061
rect 7009 24052 7021 24055
rect 6972 24024 7021 24052
rect 6972 24012 6978 24024
rect 7009 24021 7021 24024
rect 7055 24021 7067 24055
rect 7009 24015 7067 24021
rect 9030 24012 9036 24064
rect 9088 24012 9094 24064
rect 12618 24012 12624 24064
rect 12676 24012 12682 24064
rect 13751 24055 13809 24061
rect 13751 24021 13763 24055
rect 13797 24052 13809 24055
rect 13906 24052 13912 24064
rect 13797 24024 13912 24052
rect 13797 24021 13809 24024
rect 13751 24015 13809 24021
rect 13906 24012 13912 24024
rect 13964 24012 13970 24064
rect 15470 24012 15476 24064
rect 15528 24052 15534 24064
rect 17880 24052 17908 24092
rect 19150 24080 19156 24132
rect 19208 24120 19214 24132
rect 20073 24123 20131 24129
rect 20073 24120 20085 24123
rect 19208 24092 20085 24120
rect 19208 24080 19214 24092
rect 20073 24089 20085 24092
rect 20119 24089 20131 24123
rect 20272 24120 20300 24160
rect 20349 24157 20361 24191
rect 20395 24157 20407 24191
rect 20349 24151 20407 24157
rect 20438 24148 20444 24200
rect 20496 24148 20502 24200
rect 20530 24148 20536 24200
rect 20588 24148 20594 24200
rect 20809 24191 20867 24197
rect 20809 24157 20821 24191
rect 20855 24157 20867 24191
rect 20809 24151 20867 24157
rect 22097 24191 22155 24197
rect 22097 24157 22109 24191
rect 22143 24188 22155 24191
rect 22925 24191 22983 24197
rect 22143 24160 22232 24188
rect 22143 24157 22155 24160
rect 22097 24151 22155 24157
rect 20824 24120 20852 24151
rect 20272 24092 20852 24120
rect 20073 24083 20131 24089
rect 22204 24064 22232 24160
rect 22925 24157 22937 24191
rect 22971 24157 22983 24191
rect 22925 24151 22983 24157
rect 22940 24120 22968 24151
rect 23474 24148 23480 24200
rect 23532 24148 23538 24200
rect 23661 24191 23719 24197
rect 23661 24157 23673 24191
rect 23707 24188 23719 24191
rect 23750 24188 23756 24200
rect 23707 24160 23756 24188
rect 23707 24157 23719 24160
rect 23661 24151 23719 24157
rect 23750 24148 23756 24160
rect 23808 24148 23814 24200
rect 23934 24148 23940 24200
rect 23992 24148 23998 24200
rect 24210 24148 24216 24200
rect 24268 24148 24274 24200
rect 24780 24197 24808 24228
rect 25593 24225 25605 24259
rect 25639 24225 25651 24259
rect 25593 24219 25651 24225
rect 25869 24259 25927 24265
rect 25869 24225 25881 24259
rect 25915 24256 25927 24259
rect 25958 24256 25964 24268
rect 25915 24228 25964 24256
rect 25915 24225 25927 24228
rect 25869 24219 25927 24225
rect 25958 24216 25964 24228
rect 26016 24216 26022 24268
rect 26988 24256 27016 24284
rect 27338 24256 27344 24268
rect 26988 24228 27344 24256
rect 27338 24216 27344 24228
rect 27396 24216 27402 24268
rect 28261 24259 28319 24265
rect 28261 24225 28273 24259
rect 28307 24256 28319 24259
rect 28307 24228 29684 24256
rect 28307 24225 28319 24228
rect 28261 24219 28319 24225
rect 24765 24191 24823 24197
rect 24765 24157 24777 24191
rect 24811 24157 24823 24191
rect 24765 24151 24823 24157
rect 25314 24148 25320 24200
rect 25372 24148 25378 24200
rect 28166 24148 28172 24200
rect 28224 24148 28230 24200
rect 28442 24148 28448 24200
rect 28500 24148 28506 24200
rect 29454 24148 29460 24200
rect 29512 24188 29518 24200
rect 29549 24191 29607 24197
rect 29549 24188 29561 24191
rect 29512 24160 29561 24188
rect 29512 24148 29518 24160
rect 29549 24157 29561 24160
rect 29595 24157 29607 24191
rect 29656 24188 29684 24228
rect 29730 24197 29736 24200
rect 29728 24188 29736 24197
rect 29656 24160 29736 24188
rect 29549 24151 29607 24157
rect 29728 24151 29736 24160
rect 29730 24148 29736 24151
rect 29788 24148 29794 24200
rect 29840 24197 29868 24296
rect 30098 24284 30104 24296
rect 30156 24284 30162 24336
rect 31220 24324 31248 24352
rect 31772 24324 31800 24355
rect 31220 24296 31800 24324
rect 29825 24191 29883 24197
rect 29825 24157 29837 24191
rect 29871 24157 29883 24191
rect 29825 24151 29883 24157
rect 29914 24148 29920 24200
rect 29972 24148 29978 24200
rect 31404 24197 31432 24296
rect 31772 24256 31800 24296
rect 31772 24228 32444 24256
rect 32416 24197 32444 24228
rect 32785 24200 32813 24364
rect 33502 24284 33508 24336
rect 33560 24284 33566 24336
rect 34440 24333 34468 24364
rect 33689 24327 33747 24333
rect 33689 24293 33701 24327
rect 33735 24324 33747 24327
rect 34425 24327 34483 24333
rect 33735 24296 34192 24324
rect 33735 24293 33747 24296
rect 33689 24287 33747 24293
rect 33042 24216 33048 24268
rect 33100 24256 33106 24268
rect 33100 24228 34100 24256
rect 33100 24216 33106 24228
rect 31389 24191 31447 24197
rect 31389 24157 31401 24191
rect 31435 24157 31447 24191
rect 31389 24151 31447 24157
rect 31573 24191 31631 24197
rect 31573 24157 31585 24191
rect 31619 24188 31631 24191
rect 31665 24191 31723 24197
rect 31665 24188 31677 24191
rect 31619 24160 31677 24188
rect 31619 24157 31631 24160
rect 31573 24151 31631 24157
rect 31665 24157 31677 24160
rect 31711 24188 31723 24191
rect 32217 24191 32275 24197
rect 32217 24188 32229 24191
rect 31711 24160 32229 24188
rect 31711 24157 31723 24160
rect 31665 24151 31723 24157
rect 32217 24157 32229 24160
rect 32263 24157 32275 24191
rect 32217 24151 32275 24157
rect 32401 24191 32459 24197
rect 32401 24157 32413 24191
rect 32447 24157 32459 24191
rect 32401 24151 32459 24157
rect 23952 24120 23980 24148
rect 27430 24120 27436 24132
rect 22940 24092 23980 24120
rect 27094 24092 27436 24120
rect 27430 24080 27436 24092
rect 27488 24080 27494 24132
rect 31680 24120 31708 24151
rect 32766 24148 32772 24200
rect 32824 24148 32830 24200
rect 32861 24191 32919 24197
rect 32861 24157 32873 24191
rect 32907 24188 32919 24191
rect 32950 24188 32956 24200
rect 32907 24160 32956 24188
rect 32907 24157 32919 24160
rect 32861 24151 32919 24157
rect 32950 24148 32956 24160
rect 33008 24148 33014 24200
rect 33134 24148 33140 24200
rect 33192 24148 33198 24200
rect 33229 24191 33287 24197
rect 33229 24157 33241 24191
rect 33275 24157 33287 24191
rect 33229 24151 33287 24157
rect 33244 24120 33272 24151
rect 33318 24148 33324 24200
rect 33376 24188 33382 24200
rect 33597 24191 33655 24197
rect 33597 24188 33609 24191
rect 33376 24160 33609 24188
rect 33376 24148 33382 24160
rect 33597 24157 33609 24160
rect 33643 24157 33655 24191
rect 33597 24151 33655 24157
rect 33778 24148 33784 24200
rect 33836 24188 33842 24200
rect 34072 24197 34100 24228
rect 34164 24197 34192 24296
rect 34425 24293 34437 24327
rect 34471 24293 34483 24327
rect 34425 24287 34483 24293
rect 33873 24191 33931 24197
rect 33873 24188 33885 24191
rect 33836 24160 33885 24188
rect 33836 24148 33842 24160
rect 33873 24157 33885 24160
rect 33919 24157 33931 24191
rect 33873 24151 33931 24157
rect 34057 24191 34115 24197
rect 34057 24157 34069 24191
rect 34103 24157 34115 24191
rect 34057 24151 34115 24157
rect 34149 24191 34207 24197
rect 34149 24157 34161 24191
rect 34195 24157 34207 24191
rect 34149 24151 34207 24157
rect 34333 24191 34391 24197
rect 34333 24157 34345 24191
rect 34379 24157 34391 24191
rect 34333 24151 34391 24157
rect 27632 24092 31708 24120
rect 32140 24092 33272 24120
rect 33505 24123 33563 24129
rect 27632 24064 27660 24092
rect 15528 24024 17908 24052
rect 18325 24055 18383 24061
rect 15528 24012 15534 24024
rect 18325 24021 18337 24055
rect 18371 24052 18383 24055
rect 19058 24052 19064 24064
rect 18371 24024 19064 24052
rect 18371 24021 18383 24024
rect 18325 24015 18383 24021
rect 19058 24012 19064 24024
rect 19116 24012 19122 24064
rect 19242 24012 19248 24064
rect 19300 24012 19306 24064
rect 19613 24055 19671 24061
rect 19613 24021 19625 24055
rect 19659 24052 19671 24055
rect 20162 24052 20168 24064
rect 19659 24024 20168 24052
rect 19659 24021 19671 24024
rect 19613 24015 19671 24021
rect 20162 24012 20168 24024
rect 20220 24012 20226 24064
rect 22186 24012 22192 24064
rect 22244 24012 22250 24064
rect 25225 24055 25283 24061
rect 25225 24021 25237 24055
rect 25271 24052 25283 24055
rect 26510 24052 26516 24064
rect 25271 24024 26516 24052
rect 25271 24021 25283 24024
rect 25225 24015 25283 24021
rect 26510 24012 26516 24024
rect 26568 24012 26574 24064
rect 27614 24012 27620 24064
rect 27672 24012 27678 24064
rect 30190 24012 30196 24064
rect 30248 24012 30254 24064
rect 31478 24012 31484 24064
rect 31536 24012 31542 24064
rect 32140 24061 32168 24092
rect 33152 24064 33180 24092
rect 33505 24089 33517 24123
rect 33551 24120 33563 24123
rect 33965 24123 34023 24129
rect 33965 24120 33977 24123
rect 33551 24092 33977 24120
rect 33551 24089 33563 24092
rect 33505 24083 33563 24089
rect 33965 24089 33977 24092
rect 34011 24120 34023 24123
rect 34348 24120 34376 24151
rect 34011 24092 34376 24120
rect 34011 24089 34023 24092
rect 33965 24083 34023 24089
rect 32125 24055 32183 24061
rect 32125 24021 32137 24055
rect 32171 24021 32183 24055
rect 32125 24015 32183 24021
rect 32398 24012 32404 24064
rect 32456 24012 32462 24064
rect 32582 24012 32588 24064
rect 32640 24012 32646 24064
rect 33134 24012 33140 24064
rect 33192 24012 33198 24064
rect 1104 23962 38272 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38272 23962
rect 1104 23888 38272 23910
rect 1946 23808 1952 23860
rect 2004 23808 2010 23860
rect 5902 23808 5908 23860
rect 5960 23848 5966 23860
rect 6365 23851 6423 23857
rect 6365 23848 6377 23851
rect 5960 23820 6377 23848
rect 5960 23808 5966 23820
rect 6365 23817 6377 23820
rect 6411 23817 6423 23851
rect 6365 23811 6423 23817
rect 6733 23851 6791 23857
rect 6733 23817 6745 23851
rect 6779 23848 6791 23851
rect 6914 23848 6920 23860
rect 6779 23820 6920 23848
rect 6779 23817 6791 23820
rect 6733 23811 6791 23817
rect 6914 23808 6920 23820
rect 6972 23808 6978 23860
rect 7282 23808 7288 23860
rect 7340 23848 7346 23860
rect 9950 23848 9956 23860
rect 7340 23820 9956 23848
rect 7340 23808 7346 23820
rect 1964 23780 1992 23808
rect 9030 23780 9036 23792
rect 1964 23752 7604 23780
rect 5626 23672 5632 23724
rect 5684 23672 5690 23724
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23712 6883 23715
rect 7006 23712 7012 23724
rect 6871 23684 7012 23712
rect 6871 23681 6883 23684
rect 6825 23675 6883 23681
rect 7006 23672 7012 23684
rect 7064 23672 7070 23724
rect 3970 23604 3976 23656
rect 4028 23644 4034 23656
rect 6917 23647 6975 23653
rect 6917 23644 6929 23647
rect 4028 23616 6929 23644
rect 4028 23604 4034 23616
rect 6917 23613 6929 23616
rect 6963 23613 6975 23647
rect 6917 23607 6975 23613
rect 5994 23536 6000 23588
rect 6052 23576 6058 23588
rect 7282 23576 7288 23588
rect 6052 23548 7288 23576
rect 6052 23536 6058 23548
rect 7282 23536 7288 23548
rect 7340 23536 7346 23588
rect 5258 23468 5264 23520
rect 5316 23508 5322 23520
rect 5537 23511 5595 23517
rect 5537 23508 5549 23511
rect 5316 23480 5549 23508
rect 5316 23468 5322 23480
rect 5537 23477 5549 23480
rect 5583 23477 5595 23511
rect 7576 23508 7604 23752
rect 8680 23752 9036 23780
rect 8680 23721 8708 23752
rect 9030 23740 9036 23752
rect 9088 23740 9094 23792
rect 9140 23780 9168 23820
rect 9950 23808 9956 23820
rect 10008 23808 10014 23860
rect 10413 23851 10471 23857
rect 10413 23817 10425 23851
rect 10459 23848 10471 23851
rect 14737 23851 14795 23857
rect 14737 23848 14749 23851
rect 10459 23820 11192 23848
rect 10459 23817 10471 23820
rect 10413 23811 10471 23817
rect 9140 23752 9430 23780
rect 11164 23724 11192 23820
rect 13924 23820 14749 23848
rect 13924 23792 13952 23820
rect 14737 23817 14749 23820
rect 14783 23848 14795 23851
rect 14826 23848 14832 23860
rect 14783 23820 14832 23848
rect 14783 23817 14795 23820
rect 14737 23811 14795 23817
rect 14826 23808 14832 23820
rect 14884 23808 14890 23860
rect 15654 23808 15660 23860
rect 15712 23848 15718 23860
rect 15749 23851 15807 23857
rect 15749 23848 15761 23851
rect 15712 23820 15761 23848
rect 15712 23808 15718 23820
rect 15749 23817 15761 23820
rect 15795 23817 15807 23851
rect 15749 23811 15807 23817
rect 15930 23808 15936 23860
rect 15988 23848 15994 23860
rect 16942 23848 16948 23860
rect 15988 23820 16948 23848
rect 15988 23808 15994 23820
rect 16942 23808 16948 23820
rect 17000 23808 17006 23860
rect 17034 23808 17040 23860
rect 17092 23848 17098 23860
rect 17092 23820 18184 23848
rect 17092 23808 17098 23820
rect 12710 23740 12716 23792
rect 12768 23740 12774 23792
rect 13446 23740 13452 23792
rect 13504 23740 13510 23792
rect 13906 23740 13912 23792
rect 13964 23740 13970 23792
rect 14274 23740 14280 23792
rect 14332 23740 14338 23792
rect 14458 23740 14464 23792
rect 14516 23780 14522 23792
rect 14645 23783 14703 23789
rect 14645 23780 14657 23783
rect 14516 23752 14657 23780
rect 14516 23740 14522 23752
rect 14645 23749 14657 23752
rect 14691 23749 14703 23783
rect 14645 23743 14703 23749
rect 15010 23740 15016 23792
rect 15068 23740 15074 23792
rect 16025 23783 16083 23789
rect 16025 23780 16037 23783
rect 15580 23752 16037 23780
rect 8665 23715 8723 23721
rect 8665 23681 8677 23715
rect 8711 23681 8723 23715
rect 8665 23675 8723 23681
rect 11146 23672 11152 23724
rect 11204 23672 11210 23724
rect 12728 23712 12756 23740
rect 12894 23712 12900 23724
rect 12728 23684 12900 23712
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 12986 23672 12992 23724
rect 13044 23672 13050 23724
rect 14182 23672 14188 23724
rect 14240 23672 14246 23724
rect 8941 23647 8999 23653
rect 8941 23613 8953 23647
rect 8987 23644 8999 23647
rect 9306 23644 9312 23656
rect 8987 23616 9312 23644
rect 8987 23613 8999 23616
rect 8941 23607 8999 23613
rect 9306 23604 9312 23616
rect 9364 23604 9370 23656
rect 9968 23616 10732 23644
rect 9968 23508 9996 23616
rect 10042 23536 10048 23588
rect 10100 23576 10106 23588
rect 10597 23579 10655 23585
rect 10597 23576 10609 23579
rect 10100 23548 10609 23576
rect 10100 23536 10106 23548
rect 10597 23545 10609 23548
rect 10643 23545 10655 23579
rect 10597 23539 10655 23545
rect 7576 23480 9996 23508
rect 10704 23508 10732 23616
rect 12526 23604 12532 23656
rect 12584 23644 12590 23656
rect 13722 23644 13728 23656
rect 12584 23616 13728 23644
rect 12584 23604 12590 23616
rect 13722 23604 13728 23616
rect 13780 23604 13786 23656
rect 14481 23576 14509 23740
rect 14829 23715 14887 23721
rect 14829 23681 14841 23715
rect 14875 23712 14887 23715
rect 14918 23712 14924 23724
rect 14875 23684 14924 23712
rect 14875 23681 14887 23684
rect 14829 23675 14887 23681
rect 14918 23672 14924 23684
rect 14976 23672 14982 23724
rect 15102 23672 15108 23724
rect 15160 23672 15166 23724
rect 15286 23672 15292 23724
rect 15344 23672 15350 23724
rect 15470 23672 15476 23724
rect 15528 23672 15534 23724
rect 14550 23604 14556 23656
rect 14608 23644 14614 23656
rect 15120 23644 15148 23672
rect 15580 23644 15608 23752
rect 16025 23749 16037 23752
rect 16071 23780 16083 23783
rect 16850 23780 16856 23792
rect 16071 23752 16856 23780
rect 16071 23749 16083 23752
rect 16025 23743 16083 23749
rect 16850 23740 16856 23752
rect 16908 23740 16914 23792
rect 17770 23780 17776 23792
rect 17328 23752 17776 23780
rect 15657 23715 15715 23721
rect 15657 23681 15669 23715
rect 15703 23681 15715 23715
rect 15657 23675 15715 23681
rect 14608 23616 15608 23644
rect 14608 23604 14614 23616
rect 15672 23576 15700 23675
rect 16758 23672 16764 23724
rect 16816 23712 16822 23724
rect 17328 23721 17356 23752
rect 17770 23740 17776 23752
rect 17828 23740 17834 23792
rect 17313 23715 17371 23721
rect 17313 23712 17325 23715
rect 16816 23684 17325 23712
rect 16816 23672 16822 23684
rect 17313 23681 17325 23684
rect 17359 23681 17371 23715
rect 17313 23675 17371 23681
rect 17405 23715 17463 23721
rect 17405 23681 17417 23715
rect 17451 23712 17463 23715
rect 17678 23712 17684 23724
rect 17451 23684 17684 23712
rect 17451 23681 17463 23684
rect 17405 23675 17463 23681
rect 17678 23672 17684 23684
rect 17736 23712 17742 23724
rect 17957 23715 18015 23721
rect 17957 23712 17969 23715
rect 17736 23684 17969 23712
rect 17736 23672 17742 23684
rect 17957 23681 17969 23684
rect 18003 23681 18015 23715
rect 18069 23715 18127 23721
rect 18069 23712 18081 23715
rect 17957 23675 18015 23681
rect 18064 23681 18081 23712
rect 18115 23681 18127 23715
rect 18064 23675 18127 23681
rect 15841 23647 15899 23653
rect 15841 23613 15853 23647
rect 15887 23644 15899 23647
rect 16022 23644 16028 23656
rect 15887 23616 16028 23644
rect 15887 23613 15899 23616
rect 15841 23607 15899 23613
rect 16022 23604 16028 23616
rect 16080 23644 16086 23656
rect 17221 23647 17279 23653
rect 17221 23644 17233 23647
rect 16080 23616 17233 23644
rect 16080 23604 16086 23616
rect 17221 23613 17233 23616
rect 17267 23644 17279 23647
rect 17267 23616 17356 23644
rect 17267 23613 17279 23616
rect 17221 23607 17279 23613
rect 17328 23588 17356 23616
rect 17494 23604 17500 23656
rect 17552 23644 17558 23656
rect 18064 23644 18092 23675
rect 17552 23616 18092 23644
rect 18156 23644 18184 23820
rect 18690 23808 18696 23860
rect 18748 23808 18754 23860
rect 19242 23808 19248 23860
rect 19300 23808 19306 23860
rect 19334 23808 19340 23860
rect 19392 23808 19398 23860
rect 19702 23808 19708 23860
rect 19760 23848 19766 23860
rect 19981 23851 20039 23857
rect 19981 23848 19993 23851
rect 19760 23820 19993 23848
rect 19760 23808 19766 23820
rect 19981 23817 19993 23820
rect 20027 23848 20039 23851
rect 20530 23848 20536 23860
rect 20027 23820 20536 23848
rect 20027 23817 20039 23820
rect 19981 23811 20039 23817
rect 20530 23808 20536 23820
rect 20588 23808 20594 23860
rect 23106 23808 23112 23860
rect 23164 23848 23170 23860
rect 23382 23848 23388 23860
rect 23164 23820 23388 23848
rect 23164 23808 23170 23820
rect 23382 23808 23388 23820
rect 23440 23808 23446 23860
rect 23860 23820 26188 23848
rect 19260 23780 19288 23808
rect 20162 23780 20168 23792
rect 19076 23752 19288 23780
rect 19352 23752 19840 23780
rect 19076 23721 19104 23752
rect 19352 23724 19380 23752
rect 19061 23715 19119 23721
rect 19061 23681 19073 23715
rect 19107 23681 19119 23715
rect 19061 23675 19119 23681
rect 19150 23672 19156 23724
rect 19208 23672 19214 23724
rect 19334 23672 19340 23724
rect 19392 23672 19398 23724
rect 19429 23715 19487 23721
rect 19429 23681 19441 23715
rect 19475 23712 19487 23715
rect 19518 23712 19524 23724
rect 19475 23684 19524 23712
rect 19475 23681 19487 23684
rect 19429 23675 19487 23681
rect 19518 23672 19524 23684
rect 19576 23672 19582 23724
rect 19812 23721 19840 23752
rect 19904 23752 20168 23780
rect 19904 23721 19932 23752
rect 20162 23740 20168 23752
rect 20220 23740 20226 23792
rect 20254 23740 20260 23792
rect 20312 23780 20318 23792
rect 21085 23783 21143 23789
rect 20312 23752 20668 23780
rect 20312 23740 20318 23752
rect 19797 23715 19855 23721
rect 19797 23681 19809 23715
rect 19843 23681 19855 23715
rect 19797 23675 19855 23681
rect 19889 23715 19947 23721
rect 19889 23681 19901 23715
rect 19935 23681 19947 23715
rect 19889 23675 19947 23681
rect 19904 23644 19932 23675
rect 20257 23647 20315 23653
rect 20257 23644 20269 23647
rect 18156 23616 19932 23644
rect 20088 23616 20269 23644
rect 17552 23604 17558 23616
rect 14481 23548 16436 23576
rect 12713 23511 12771 23517
rect 12713 23508 12725 23511
rect 10704 23480 12725 23508
rect 5537 23471 5595 23477
rect 12713 23477 12725 23480
rect 12759 23477 12771 23511
rect 12713 23471 12771 23477
rect 14826 23468 14832 23520
rect 14884 23508 14890 23520
rect 15105 23511 15163 23517
rect 15105 23508 15117 23511
rect 14884 23480 15117 23508
rect 14884 23468 14890 23480
rect 15105 23477 15117 23480
rect 15151 23477 15163 23511
rect 15105 23471 15163 23477
rect 15933 23511 15991 23517
rect 15933 23477 15945 23511
rect 15979 23508 15991 23511
rect 16206 23508 16212 23520
rect 15979 23480 16212 23508
rect 15979 23477 15991 23480
rect 15933 23471 15991 23477
rect 16206 23468 16212 23480
rect 16264 23468 16270 23520
rect 16408 23508 16436 23548
rect 17310 23536 17316 23588
rect 17368 23536 17374 23588
rect 18414 23576 18420 23588
rect 17511 23548 18420 23576
rect 17511 23508 17539 23548
rect 16408 23480 17539 23508
rect 17586 23468 17592 23520
rect 17644 23508 17650 23520
rect 17681 23511 17739 23517
rect 17681 23508 17693 23511
rect 17644 23480 17693 23508
rect 17644 23468 17650 23480
rect 17681 23477 17693 23480
rect 17727 23477 17739 23511
rect 17681 23471 17739 23477
rect 17770 23468 17776 23520
rect 17828 23468 17834 23520
rect 18248 23517 18276 23548
rect 18414 23536 18420 23548
rect 18472 23536 18478 23588
rect 18969 23579 19027 23585
rect 18969 23545 18981 23579
rect 19015 23576 19027 23579
rect 19521 23579 19579 23585
rect 19521 23576 19533 23579
rect 19015 23548 19533 23576
rect 19015 23545 19027 23548
rect 18969 23539 19027 23545
rect 19521 23545 19533 23548
rect 19567 23545 19579 23579
rect 19521 23539 19579 23545
rect 19886 23536 19892 23588
rect 19944 23576 19950 23588
rect 20088 23576 20116 23616
rect 20257 23613 20269 23616
rect 20303 23613 20315 23647
rect 20640 23644 20668 23752
rect 21085 23749 21097 23783
rect 21131 23780 21143 23783
rect 21358 23780 21364 23792
rect 21131 23752 21364 23780
rect 21131 23749 21143 23752
rect 21085 23743 21143 23749
rect 21358 23740 21364 23752
rect 21416 23740 21422 23792
rect 22373 23783 22431 23789
rect 22373 23749 22385 23783
rect 22419 23780 22431 23783
rect 22646 23780 22652 23792
rect 22419 23752 22652 23780
rect 22419 23749 22431 23752
rect 22373 23743 22431 23749
rect 22646 23740 22652 23752
rect 22704 23740 22710 23792
rect 23860 23724 23888 23820
rect 25314 23780 25320 23792
rect 24688 23752 25320 23780
rect 20806 23672 20812 23724
rect 20864 23672 20870 23724
rect 22557 23715 22615 23721
rect 22557 23681 22569 23715
rect 22603 23712 22615 23715
rect 22922 23712 22928 23724
rect 22603 23684 22928 23712
rect 22603 23681 22615 23684
rect 22557 23675 22615 23681
rect 22922 23672 22928 23684
rect 22980 23672 22986 23724
rect 23014 23672 23020 23724
rect 23072 23712 23078 23724
rect 23293 23715 23351 23721
rect 23293 23712 23305 23715
rect 23072 23684 23305 23712
rect 23072 23672 23078 23684
rect 23293 23681 23305 23684
rect 23339 23681 23351 23715
rect 23293 23675 23351 23681
rect 23661 23715 23719 23721
rect 23661 23681 23673 23715
rect 23707 23712 23719 23715
rect 23750 23712 23756 23724
rect 23707 23684 23756 23712
rect 23707 23681 23719 23684
rect 23661 23675 23719 23681
rect 23750 23672 23756 23684
rect 23808 23672 23814 23724
rect 23842 23672 23848 23724
rect 23900 23672 23906 23724
rect 24688 23721 24716 23752
rect 25314 23740 25320 23752
rect 25372 23780 25378 23792
rect 25869 23783 25927 23789
rect 25869 23780 25881 23783
rect 25372 23752 25881 23780
rect 25372 23740 25378 23752
rect 25869 23749 25881 23752
rect 25915 23749 25927 23783
rect 25869 23743 25927 23749
rect 24673 23715 24731 23721
rect 24673 23681 24685 23715
rect 24719 23681 24731 23715
rect 24673 23675 24731 23681
rect 24762 23672 24768 23724
rect 24820 23712 24826 23724
rect 25041 23715 25099 23721
rect 25041 23712 25053 23715
rect 24820 23684 25053 23712
rect 24820 23672 24826 23684
rect 25041 23681 25053 23684
rect 25087 23681 25099 23715
rect 25041 23675 25099 23681
rect 25130 23672 25136 23724
rect 25188 23672 25194 23724
rect 26050 23672 26056 23724
rect 26108 23672 26114 23724
rect 26160 23721 26188 23820
rect 26418 23808 26424 23860
rect 26476 23848 26482 23860
rect 28629 23851 28687 23857
rect 28629 23848 28641 23851
rect 26476 23820 28641 23848
rect 26476 23808 26482 23820
rect 28629 23817 28641 23820
rect 28675 23817 28687 23851
rect 28629 23811 28687 23817
rect 28810 23808 28816 23860
rect 28868 23848 28874 23860
rect 29089 23851 29147 23857
rect 29089 23848 29101 23851
rect 28868 23820 29101 23848
rect 28868 23808 28874 23820
rect 29089 23817 29101 23820
rect 29135 23817 29147 23851
rect 29089 23811 29147 23817
rect 31478 23808 31484 23860
rect 31536 23848 31542 23860
rect 32217 23851 32275 23857
rect 31536 23820 31754 23848
rect 31536 23808 31542 23820
rect 27154 23780 27160 23792
rect 26252 23752 27160 23780
rect 26145 23715 26203 23721
rect 26145 23681 26157 23715
rect 26191 23681 26203 23715
rect 26145 23675 26203 23681
rect 24400 23656 24452 23662
rect 22649 23647 22707 23653
rect 22649 23644 22661 23647
rect 20640 23616 22661 23644
rect 20257 23607 20315 23613
rect 22649 23613 22661 23616
rect 22695 23613 22707 23647
rect 22649 23607 22707 23613
rect 23201 23647 23259 23653
rect 23201 23613 23213 23647
rect 23247 23613 23259 23647
rect 23201 23607 23259 23613
rect 19944 23548 20116 23576
rect 20165 23579 20223 23585
rect 19944 23536 19950 23548
rect 20165 23545 20177 23579
rect 20211 23576 20223 23579
rect 20346 23576 20352 23588
rect 20211 23548 20352 23576
rect 20211 23545 20223 23548
rect 20165 23539 20223 23545
rect 20346 23536 20352 23548
rect 20404 23536 20410 23588
rect 22186 23536 22192 23588
rect 22244 23576 22250 23588
rect 23216 23576 23244 23607
rect 25866 23604 25872 23656
rect 25924 23644 25930 23656
rect 26252 23644 26280 23752
rect 27154 23740 27160 23752
rect 27212 23780 27218 23792
rect 27249 23783 27307 23789
rect 27249 23780 27261 23783
rect 27212 23752 27261 23780
rect 27212 23740 27218 23752
rect 27249 23749 27261 23752
rect 27295 23749 27307 23783
rect 28166 23780 28172 23792
rect 27249 23743 27307 23749
rect 27540 23752 28172 23780
rect 27540 23724 27568 23752
rect 27062 23672 27068 23724
rect 27120 23672 27126 23724
rect 27341 23715 27399 23721
rect 27341 23712 27353 23715
rect 27172 23684 27353 23712
rect 27172 23644 27200 23684
rect 27341 23681 27353 23684
rect 27387 23681 27399 23715
rect 27341 23675 27399 23681
rect 27433 23715 27491 23721
rect 27433 23681 27445 23715
rect 27479 23712 27491 23715
rect 27522 23712 27528 23724
rect 27479 23684 27528 23712
rect 27479 23681 27491 23684
rect 27433 23675 27491 23681
rect 27522 23672 27528 23684
rect 27580 23672 27586 23724
rect 27706 23672 27712 23724
rect 27764 23672 27770 23724
rect 28092 23721 28120 23752
rect 28166 23740 28172 23752
rect 28224 23740 28230 23792
rect 28721 23783 28779 23789
rect 28721 23749 28733 23783
rect 28767 23780 28779 23783
rect 28902 23780 28908 23792
rect 28767 23752 28908 23780
rect 28767 23749 28779 23752
rect 28721 23743 28779 23749
rect 28902 23740 28908 23752
rect 28960 23740 28966 23792
rect 27893 23715 27951 23721
rect 27893 23681 27905 23715
rect 27939 23681 27951 23715
rect 27893 23675 27951 23681
rect 27985 23715 28043 23721
rect 27985 23681 27997 23715
rect 28031 23681 28043 23715
rect 27985 23675 28043 23681
rect 28077 23715 28135 23721
rect 28077 23681 28089 23715
rect 28123 23681 28135 23715
rect 31726 23712 31754 23820
rect 32217 23817 32229 23851
rect 32263 23848 32275 23851
rect 32950 23848 32956 23860
rect 32263 23820 32956 23848
rect 32263 23817 32275 23820
rect 32217 23811 32275 23817
rect 32950 23808 32956 23820
rect 33008 23808 33014 23860
rect 33134 23808 33140 23860
rect 33192 23808 33198 23860
rect 33152 23721 33180 23808
rect 32125 23715 32183 23721
rect 32125 23712 32137 23715
rect 31726 23684 32137 23712
rect 28077 23675 28135 23681
rect 32125 23681 32137 23684
rect 32171 23681 32183 23715
rect 32125 23675 32183 23681
rect 33137 23715 33195 23721
rect 33137 23681 33149 23715
rect 33183 23681 33195 23715
rect 33137 23675 33195 23681
rect 27908 23644 27936 23675
rect 25924 23616 26280 23644
rect 26344 23616 27200 23644
rect 27356 23616 27936 23644
rect 25924 23604 25930 23616
rect 24400 23598 24452 23604
rect 22244 23548 23244 23576
rect 22244 23536 22250 23548
rect 24302 23536 24308 23588
rect 24360 23536 24366 23588
rect 18233 23511 18291 23517
rect 18233 23477 18245 23511
rect 18279 23477 18291 23511
rect 18233 23471 18291 23477
rect 19794 23468 19800 23520
rect 19852 23508 19858 23520
rect 26344 23508 26372 23616
rect 27154 23536 27160 23588
rect 27212 23576 27218 23588
rect 27356 23576 27384 23616
rect 27212 23548 27384 23576
rect 27212 23536 27218 23548
rect 27430 23536 27436 23588
rect 27488 23536 27494 23588
rect 27614 23536 27620 23588
rect 27672 23536 27678 23588
rect 27706 23536 27712 23588
rect 27764 23576 27770 23588
rect 28000 23576 28028 23675
rect 34606 23672 34612 23724
rect 34664 23712 34670 23724
rect 35529 23715 35587 23721
rect 35529 23712 35541 23715
rect 34664 23684 35541 23712
rect 34664 23672 34670 23684
rect 35529 23681 35541 23684
rect 35575 23681 35587 23715
rect 35529 23675 35587 23681
rect 28445 23647 28503 23653
rect 28445 23644 28457 23647
rect 27764 23548 28028 23576
rect 28184 23616 28457 23644
rect 27764 23536 27770 23548
rect 19852 23480 26372 23508
rect 27448 23508 27476 23536
rect 28184 23508 28212 23616
rect 28445 23613 28457 23616
rect 28491 23644 28503 23647
rect 33410 23644 33416 23656
rect 28491 23616 33416 23644
rect 28491 23613 28503 23616
rect 28445 23607 28503 23613
rect 33410 23604 33416 23616
rect 33468 23604 33474 23656
rect 34977 23647 35035 23653
rect 34977 23613 34989 23647
rect 35023 23644 35035 23647
rect 35342 23644 35348 23656
rect 35023 23616 35348 23644
rect 35023 23613 35035 23616
rect 34977 23607 35035 23613
rect 35342 23604 35348 23616
rect 35400 23604 35406 23656
rect 35802 23604 35808 23656
rect 35860 23604 35866 23656
rect 28261 23579 28319 23585
rect 28261 23545 28273 23579
rect 28307 23576 28319 23579
rect 33042 23576 33048 23588
rect 28307 23548 33048 23576
rect 28307 23545 28319 23548
rect 28261 23539 28319 23545
rect 33042 23536 33048 23548
rect 33100 23536 33106 23588
rect 27448 23480 28212 23508
rect 19852 23468 19858 23480
rect 33226 23468 33232 23520
rect 33284 23468 33290 23520
rect 1104 23418 38272 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38272 23418
rect 1104 23344 38272 23366
rect 1762 23264 1768 23316
rect 1820 23304 1826 23316
rect 2225 23307 2283 23313
rect 2225 23304 2237 23307
rect 1820 23276 2237 23304
rect 1820 23264 1826 23276
rect 2225 23273 2237 23276
rect 2271 23273 2283 23307
rect 2225 23267 2283 23273
rect 2774 23264 2780 23316
rect 2832 23304 2838 23316
rect 2961 23307 3019 23313
rect 2961 23304 2973 23307
rect 2832 23276 2973 23304
rect 2832 23264 2838 23276
rect 2961 23273 2973 23276
rect 3007 23273 3019 23307
rect 4154 23304 4160 23316
rect 2961 23267 3019 23273
rect 3068 23276 4160 23304
rect 1946 23060 1952 23112
rect 2004 23060 2010 23112
rect 2501 23103 2559 23109
rect 2501 23069 2513 23103
rect 2547 23069 2559 23103
rect 2501 23063 2559 23069
rect 2593 23103 2651 23109
rect 2593 23069 2605 23103
rect 2639 23069 2651 23103
rect 2593 23063 2651 23069
rect 2516 22976 2544 23063
rect 2608 23032 2636 23063
rect 2682 23060 2688 23112
rect 2740 23060 2746 23112
rect 2869 23103 2927 23109
rect 2869 23069 2881 23103
rect 2915 23100 2927 23103
rect 3068 23100 3096 23276
rect 4154 23264 4160 23276
rect 4212 23264 4218 23316
rect 4249 23307 4307 23313
rect 4249 23273 4261 23307
rect 4295 23304 4307 23307
rect 4614 23304 4620 23316
rect 4295 23276 4620 23304
rect 4295 23273 4307 23276
rect 4249 23267 4307 23273
rect 4614 23264 4620 23276
rect 4672 23264 4678 23316
rect 4798 23264 4804 23316
rect 4856 23304 4862 23316
rect 4985 23307 5043 23313
rect 4985 23304 4997 23307
rect 4856 23276 4997 23304
rect 4856 23264 4862 23276
rect 4985 23273 4997 23276
rect 5031 23273 5043 23307
rect 4985 23267 5043 23273
rect 5626 23264 5632 23316
rect 5684 23304 5690 23316
rect 6273 23307 6331 23313
rect 6273 23304 6285 23307
rect 5684 23276 6285 23304
rect 5684 23264 5690 23276
rect 6273 23273 6285 23276
rect 6319 23273 6331 23307
rect 6457 23307 6515 23313
rect 6457 23304 6469 23307
rect 6273 23267 6331 23273
rect 6380 23276 6469 23304
rect 5350 23236 5356 23248
rect 3344 23208 5356 23236
rect 2915 23072 3096 23100
rect 2915 23069 2927 23072
rect 2869 23063 2927 23069
rect 3142 23060 3148 23112
rect 3200 23060 3206 23112
rect 3344 23109 3372 23208
rect 3329 23103 3387 23109
rect 3329 23069 3341 23103
rect 3375 23069 3387 23103
rect 3329 23063 3387 23069
rect 3602 23060 3608 23112
rect 3660 23060 3666 23112
rect 4430 23060 4436 23112
rect 4488 23060 4494 23112
rect 4632 23109 4660 23208
rect 5350 23196 5356 23208
rect 5408 23196 5414 23248
rect 5810 23196 5816 23248
rect 5868 23236 5874 23248
rect 6380 23236 6408 23276
rect 6457 23273 6469 23276
rect 6503 23273 6515 23307
rect 6457 23267 6515 23273
rect 7006 23264 7012 23316
rect 7064 23264 7070 23316
rect 7190 23264 7196 23316
rect 7248 23304 7254 23316
rect 8113 23307 8171 23313
rect 8113 23304 8125 23307
rect 7248 23276 8125 23304
rect 7248 23264 7254 23276
rect 8113 23273 8125 23276
rect 8159 23273 8171 23307
rect 8113 23267 8171 23273
rect 9306 23264 9312 23316
rect 9364 23264 9370 23316
rect 9398 23264 9404 23316
rect 9456 23304 9462 23316
rect 14093 23307 14151 23313
rect 9456 23276 14044 23304
rect 9456 23264 9462 23276
rect 5868 23208 6408 23236
rect 6748 23208 7696 23236
rect 5868 23196 5874 23208
rect 5721 23171 5779 23177
rect 5721 23168 5733 23171
rect 5184 23140 5733 23168
rect 4617 23103 4675 23109
rect 4617 23069 4629 23103
rect 4663 23069 4675 23103
rect 4617 23063 4675 23069
rect 4890 23060 4896 23112
rect 4948 23060 4954 23112
rect 5184 23109 5212 23140
rect 5721 23137 5733 23140
rect 5767 23137 5779 23171
rect 6546 23168 6552 23180
rect 5721 23131 5779 23137
rect 5828 23140 6552 23168
rect 5169 23103 5227 23109
rect 5169 23069 5181 23103
rect 5215 23069 5227 23103
rect 5169 23063 5227 23069
rect 5629 23103 5687 23109
rect 5629 23069 5641 23103
rect 5675 23100 5687 23103
rect 5828 23100 5856 23140
rect 6546 23128 6552 23140
rect 6604 23128 6610 23180
rect 5675 23072 5856 23100
rect 5675 23069 5687 23072
rect 5629 23063 5687 23069
rect 5902 23060 5908 23112
rect 5960 23060 5966 23112
rect 6748 23109 6776 23208
rect 7668 23168 7696 23208
rect 10134 23196 10140 23248
rect 10192 23236 10198 23248
rect 10594 23236 10600 23248
rect 10192 23208 10600 23236
rect 10192 23196 10198 23208
rect 10594 23196 10600 23208
rect 10652 23196 10658 23248
rect 14016 23236 14044 23276
rect 14093 23273 14105 23307
rect 14139 23304 14151 23307
rect 14182 23304 14188 23316
rect 14139 23276 14188 23304
rect 14139 23273 14151 23276
rect 14093 23267 14151 23273
rect 14182 23264 14188 23276
rect 14240 23264 14246 23316
rect 15010 23264 15016 23316
rect 15068 23304 15074 23316
rect 15286 23304 15292 23316
rect 15068 23276 15292 23304
rect 15068 23264 15074 23276
rect 15286 23264 15292 23276
rect 15344 23304 15350 23316
rect 16022 23304 16028 23316
rect 15344 23276 16028 23304
rect 15344 23264 15350 23276
rect 16022 23264 16028 23276
rect 16080 23264 16086 23316
rect 19794 23304 19800 23316
rect 18340 23276 19800 23304
rect 18340 23236 18368 23276
rect 19794 23264 19800 23276
rect 19852 23264 19858 23316
rect 19886 23264 19892 23316
rect 19944 23304 19950 23316
rect 20441 23307 20499 23313
rect 20441 23304 20453 23307
rect 19944 23276 20453 23304
rect 19944 23264 19950 23276
rect 20441 23273 20453 23276
rect 20487 23273 20499 23307
rect 20441 23267 20499 23273
rect 20806 23264 20812 23316
rect 20864 23264 20870 23316
rect 22554 23304 22560 23316
rect 22020 23276 22560 23304
rect 14016 23208 18368 23236
rect 7668 23140 7788 23168
rect 6181 23103 6239 23109
rect 6181 23100 6193 23103
rect 6012 23072 6193 23100
rect 3237 23035 3295 23041
rect 2608 23004 2774 23032
rect 1765 22967 1823 22973
rect 1765 22933 1777 22967
rect 1811 22964 1823 22967
rect 1854 22964 1860 22976
rect 1811 22936 1860 22964
rect 1811 22933 1823 22936
rect 1765 22927 1823 22933
rect 1854 22924 1860 22936
rect 1912 22924 1918 22976
rect 2498 22924 2504 22976
rect 2556 22924 2562 22976
rect 2746 22964 2774 23004
rect 3237 23001 3249 23035
rect 3283 23001 3295 23035
rect 3237 22995 3295 23001
rect 3467 23035 3525 23041
rect 3467 23001 3479 23035
rect 3513 23032 3525 23035
rect 3513 23004 4292 23032
rect 3513 23001 3525 23004
rect 3467 22995 3525 23001
rect 2866 22964 2872 22976
rect 2746 22936 2872 22964
rect 2866 22924 2872 22936
rect 2924 22924 2930 22976
rect 3252 22964 3280 22995
rect 3970 22964 3976 22976
rect 3252 22936 3976 22964
rect 3970 22924 3976 22936
rect 4028 22924 4034 22976
rect 4264 22964 4292 23004
rect 4522 22992 4528 23044
rect 4580 22992 4586 23044
rect 4735 23035 4793 23041
rect 4735 23032 4747 23035
rect 4632 23004 4747 23032
rect 4632 22976 4660 23004
rect 4735 23001 4747 23004
rect 4781 23001 4793 23035
rect 4735 22995 4793 23001
rect 5258 22992 5264 23044
rect 5316 22992 5322 23044
rect 5350 22992 5356 23044
rect 5408 22992 5414 23044
rect 5471 23035 5529 23041
rect 5471 23001 5483 23035
rect 5517 23001 5529 23035
rect 5471 22995 5529 23001
rect 6012 23032 6040 23072
rect 6181 23069 6193 23072
rect 6227 23069 6239 23103
rect 6733 23103 6791 23109
rect 6733 23100 6745 23103
rect 6181 23063 6239 23069
rect 6564 23072 6745 23100
rect 6425 23035 6483 23041
rect 6425 23032 6437 23035
rect 6012 23004 6437 23032
rect 4614 22964 4620 22976
rect 4264 22936 4620 22964
rect 4614 22924 4620 22936
rect 4672 22964 4678 22976
rect 5486 22964 5514 22995
rect 6012 22976 6040 23004
rect 6425 23001 6437 23004
rect 6471 23032 6483 23035
rect 6564 23032 6592 23072
rect 6733 23069 6745 23072
rect 6779 23069 6791 23103
rect 6917 23103 6975 23109
rect 6917 23100 6929 23103
rect 6733 23063 6791 23069
rect 6840 23072 6929 23100
rect 6471 23004 6592 23032
rect 6641 23035 6699 23041
rect 6471 23001 6483 23004
rect 6425 22995 6483 23001
rect 6641 23001 6653 23035
rect 6687 23032 6699 23035
rect 6840 23032 6868 23072
rect 6917 23069 6929 23072
rect 6963 23100 6975 23103
rect 7006 23100 7012 23112
rect 6963 23072 7012 23100
rect 6963 23069 6975 23072
rect 6917 23063 6975 23069
rect 7006 23060 7012 23072
rect 7064 23060 7070 23112
rect 7760 23109 7788 23140
rect 9122 23128 9128 23180
rect 9180 23168 9186 23180
rect 9180 23140 10548 23168
rect 9180 23128 9186 23140
rect 7653 23103 7711 23109
rect 7194 23081 7252 23087
rect 7194 23047 7206 23081
rect 7240 23047 7252 23081
rect 7653 23069 7665 23103
rect 7699 23069 7711 23103
rect 7653 23063 7711 23069
rect 7745 23103 7803 23109
rect 7745 23069 7757 23103
rect 7791 23069 7803 23103
rect 9398 23100 9404 23112
rect 7745 23063 7803 23069
rect 7852 23072 9404 23100
rect 7194 23044 7252 23047
rect 6687 23004 6868 23032
rect 6687 23001 6699 23004
rect 6641 22995 6699 23001
rect 4672 22936 5514 22964
rect 4672 22924 4678 22936
rect 5994 22924 6000 22976
rect 6052 22924 6058 22976
rect 6089 22967 6147 22973
rect 6089 22933 6101 22967
rect 6135 22964 6147 22967
rect 6656 22964 6684 22995
rect 7190 22992 7196 23044
rect 7248 22992 7254 23044
rect 7285 23035 7343 23041
rect 7285 23001 7297 23035
rect 7331 23001 7343 23035
rect 7285 22995 7343 23001
rect 6135 22936 6684 22964
rect 6917 22967 6975 22973
rect 6135 22933 6147 22936
rect 6089 22927 6147 22933
rect 6917 22933 6929 22967
rect 6963 22964 6975 22967
rect 7300 22964 7328 22995
rect 7374 22992 7380 23044
rect 7432 22992 7438 23044
rect 7558 23041 7564 23044
rect 7515 23035 7564 23041
rect 7515 23001 7527 23035
rect 7561 23001 7564 23035
rect 7515 22995 7564 23001
rect 7558 22992 7564 22995
rect 7616 22992 7622 23044
rect 7668 23032 7696 23063
rect 7852 23032 7880 23072
rect 9398 23060 9404 23072
rect 9456 23060 9462 23112
rect 9490 23060 9496 23112
rect 9548 23060 9554 23112
rect 9585 23103 9643 23109
rect 9585 23069 9597 23103
rect 9631 23100 9643 23103
rect 9631 23072 9812 23100
rect 9631 23069 9643 23072
rect 9585 23063 9643 23069
rect 7668 23004 7880 23032
rect 7926 22992 7932 23044
rect 7984 22992 7990 23044
rect 9674 22992 9680 23044
rect 9732 22992 9738 23044
rect 9784 23032 9812 23072
rect 9858 23060 9864 23112
rect 9916 23060 9922 23112
rect 10042 23060 10048 23112
rect 10100 23060 10106 23112
rect 10520 23109 10548 23140
rect 11146 23128 11152 23180
rect 11204 23168 11210 23180
rect 12066 23168 12072 23180
rect 11204 23140 12072 23168
rect 11204 23128 11210 23140
rect 12066 23128 12072 23140
rect 12124 23128 12130 23180
rect 12342 23128 12348 23180
rect 12400 23168 12406 23180
rect 12805 23171 12863 23177
rect 12805 23168 12817 23171
rect 12400 23140 12817 23168
rect 12400 23128 12406 23140
rect 12805 23137 12817 23140
rect 12851 23168 12863 23171
rect 15562 23168 15568 23180
rect 12851 23140 15568 23168
rect 12851 23137 12863 23140
rect 12805 23131 12863 23137
rect 15562 23128 15568 23140
rect 15620 23128 15626 23180
rect 15654 23128 15660 23180
rect 15712 23128 15718 23180
rect 16114 23128 16120 23180
rect 16172 23168 16178 23180
rect 16209 23171 16267 23177
rect 16209 23168 16221 23171
rect 16172 23140 16221 23168
rect 16172 23128 16178 23140
rect 16209 23137 16221 23140
rect 16255 23137 16267 23171
rect 16209 23131 16267 23137
rect 16684 23140 17908 23168
rect 10505 23103 10563 23109
rect 10505 23069 10517 23103
rect 10551 23069 10563 23103
rect 10505 23063 10563 23069
rect 10597 23103 10655 23109
rect 10597 23069 10609 23103
rect 10643 23100 10655 23103
rect 10781 23103 10839 23109
rect 10781 23100 10793 23103
rect 10643 23072 10793 23100
rect 10643 23069 10655 23072
rect 10597 23063 10655 23069
rect 10781 23069 10793 23072
rect 10827 23069 10839 23103
rect 10781 23063 10839 23069
rect 12710 23060 12716 23112
rect 12768 23100 12774 23112
rect 15010 23100 15016 23112
rect 12768 23072 15016 23100
rect 12768 23060 12774 23072
rect 15010 23060 15016 23072
rect 15068 23060 15074 23112
rect 15102 23060 15108 23112
rect 15160 23100 15166 23112
rect 15197 23103 15255 23109
rect 15197 23100 15209 23103
rect 15160 23072 15209 23100
rect 15160 23060 15166 23072
rect 15197 23069 15209 23072
rect 15243 23069 15255 23103
rect 15197 23063 15255 23069
rect 15378 23060 15384 23112
rect 15436 23060 15442 23112
rect 15749 23103 15807 23109
rect 15749 23100 15761 23103
rect 15488 23072 15761 23100
rect 10060 23032 10088 23060
rect 9784 23004 10088 23032
rect 11054 22992 11060 23044
rect 11112 22992 11118 23044
rect 11146 22992 11152 23044
rect 11204 23032 11210 23044
rect 11204 23004 11546 23032
rect 11204 22992 11210 23004
rect 13998 22992 14004 23044
rect 14056 23032 14062 23044
rect 14277 23035 14335 23041
rect 14277 23032 14289 23035
rect 14056 23004 14289 23032
rect 14056 22992 14062 23004
rect 14277 23001 14289 23004
rect 14323 23001 14335 23035
rect 14277 22995 14335 23001
rect 14458 22992 14464 23044
rect 14516 22992 14522 23044
rect 14642 22992 14648 23044
rect 14700 23032 14706 23044
rect 14737 23035 14795 23041
rect 14737 23032 14749 23035
rect 14700 23004 14749 23032
rect 14700 22992 14706 23004
rect 14737 23001 14749 23004
rect 14783 23001 14795 23035
rect 14737 22995 14795 23001
rect 6963 22936 7328 22964
rect 6963 22933 6975 22936
rect 6917 22927 6975 22933
rect 7650 22924 7656 22976
rect 7708 22964 7714 22976
rect 12526 22964 12532 22976
rect 7708 22936 12532 22964
rect 7708 22924 7714 22936
rect 12526 22924 12532 22936
rect 12584 22924 12590 22976
rect 13446 22924 13452 22976
rect 13504 22964 13510 22976
rect 15488 22964 15516 23072
rect 15749 23069 15761 23072
rect 15795 23100 15807 23103
rect 15838 23100 15844 23112
rect 15795 23072 15844 23100
rect 15795 23069 15807 23072
rect 15749 23063 15807 23069
rect 15838 23060 15844 23072
rect 15896 23060 15902 23112
rect 16684 23109 16712 23140
rect 17880 23112 17908 23140
rect 17954 23128 17960 23180
rect 18012 23168 18018 23180
rect 18693 23171 18751 23177
rect 18693 23168 18705 23171
rect 18012 23140 18705 23168
rect 18012 23128 18018 23140
rect 16669 23103 16727 23109
rect 16669 23069 16681 23103
rect 16715 23069 16727 23103
rect 16669 23063 16727 23069
rect 17037 23103 17095 23109
rect 17037 23069 17049 23103
rect 17083 23069 17095 23103
rect 17037 23063 17095 23069
rect 17052 23032 17080 23063
rect 17126 23060 17132 23112
rect 17184 23060 17190 23112
rect 17402 23060 17408 23112
rect 17460 23060 17466 23112
rect 17678 23060 17684 23112
rect 17736 23060 17742 23112
rect 17862 23060 17868 23112
rect 17920 23060 17926 23112
rect 18233 23103 18291 23109
rect 18233 23069 18245 23103
rect 18279 23069 18291 23103
rect 18233 23063 18291 23069
rect 17310 23032 17316 23044
rect 17052 23004 17316 23032
rect 17310 22992 17316 23004
rect 17368 22992 17374 23044
rect 17770 22992 17776 23044
rect 17828 23032 17834 23044
rect 18248 23032 18276 23063
rect 17828 23004 18276 23032
rect 18524 23032 18552 23140
rect 18693 23137 18705 23140
rect 18739 23137 18751 23171
rect 18693 23131 18751 23137
rect 20530 23128 20536 23180
rect 20588 23128 20594 23180
rect 22020 23177 22048 23276
rect 22554 23264 22560 23276
rect 22612 23304 22618 23316
rect 23290 23304 23296 23316
rect 22612 23276 23296 23304
rect 22612 23264 22618 23276
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 23382 23264 23388 23316
rect 23440 23304 23446 23316
rect 23845 23307 23903 23313
rect 23845 23304 23857 23307
rect 23440 23276 23857 23304
rect 23440 23264 23446 23276
rect 23845 23273 23857 23276
rect 23891 23304 23903 23307
rect 26050 23304 26056 23316
rect 23891 23276 26056 23304
rect 23891 23273 23903 23276
rect 23845 23267 23903 23273
rect 26050 23264 26056 23276
rect 26108 23264 26114 23316
rect 26326 23264 26332 23316
rect 26384 23304 26390 23316
rect 29362 23304 29368 23316
rect 26384 23276 29368 23304
rect 26384 23264 26390 23276
rect 29362 23264 29368 23276
rect 29420 23264 29426 23316
rect 32030 23264 32036 23316
rect 32088 23304 32094 23316
rect 33042 23304 33048 23316
rect 32088 23276 33048 23304
rect 32088 23264 32094 23276
rect 33042 23264 33048 23276
rect 33100 23264 33106 23316
rect 34606 23264 34612 23316
rect 34664 23304 34670 23316
rect 34793 23307 34851 23313
rect 34664 23276 34744 23304
rect 34664 23264 34670 23276
rect 23474 23196 23480 23248
rect 23532 23196 23538 23248
rect 27522 23196 27528 23248
rect 27580 23236 27586 23248
rect 27580 23208 34652 23236
rect 27580 23196 27586 23208
rect 22005 23171 22063 23177
rect 22005 23137 22017 23171
rect 22051 23137 22063 23171
rect 22005 23131 22063 23137
rect 22186 23128 22192 23180
rect 22244 23168 22250 23180
rect 22741 23171 22799 23177
rect 22741 23168 22753 23171
rect 22244 23140 22753 23168
rect 22244 23128 22250 23140
rect 22741 23137 22753 23140
rect 22787 23168 22799 23171
rect 23842 23168 23848 23180
rect 22787 23140 23848 23168
rect 22787 23137 22799 23140
rect 22741 23131 22799 23137
rect 23842 23128 23848 23140
rect 23900 23128 23906 23180
rect 24854 23128 24860 23180
rect 24912 23168 24918 23180
rect 24912 23140 25728 23168
rect 24912 23128 24918 23140
rect 18598 23060 18604 23112
rect 18656 23100 18662 23112
rect 20438 23100 20444 23112
rect 18656 23072 20444 23100
rect 18656 23060 18662 23072
rect 20438 23060 20444 23072
rect 20496 23060 20502 23112
rect 20622 23060 20628 23112
rect 20680 23100 20686 23112
rect 21177 23103 21235 23109
rect 21177 23100 21189 23103
rect 20680 23072 21189 23100
rect 20680 23060 20686 23072
rect 21177 23069 21189 23072
rect 21223 23069 21235 23103
rect 21177 23063 21235 23069
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23100 21787 23103
rect 22278 23100 22284 23112
rect 21775 23072 22284 23100
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 22278 23060 22284 23072
rect 22336 23060 22342 23112
rect 22922 23060 22928 23112
rect 22980 23060 22986 23112
rect 23014 23060 23020 23112
rect 23072 23100 23078 23112
rect 23385 23103 23443 23109
rect 23385 23100 23397 23103
rect 23072 23072 23397 23100
rect 23072 23060 23078 23072
rect 23385 23069 23397 23072
rect 23431 23069 23443 23103
rect 23385 23063 23443 23069
rect 23753 23103 23811 23109
rect 23753 23069 23765 23103
rect 23799 23069 23811 23103
rect 23753 23063 23811 23069
rect 23937 23103 23995 23109
rect 23937 23069 23949 23103
rect 23983 23069 23995 23103
rect 23937 23063 23995 23069
rect 19702 23032 19708 23044
rect 18524 23004 19708 23032
rect 17828 22992 17834 23004
rect 13504 22936 15516 22964
rect 13504 22924 13510 22936
rect 15562 22924 15568 22976
rect 15620 22964 15626 22976
rect 17494 22964 17500 22976
rect 15620 22936 17500 22964
rect 15620 22924 15626 22936
rect 17494 22924 17500 22936
rect 17552 22924 17558 22976
rect 18248 22964 18276 23004
rect 19702 22992 19708 23004
rect 19760 22992 19766 23044
rect 20254 22992 20260 23044
rect 20312 23032 20318 23044
rect 20993 23035 21051 23041
rect 20993 23032 21005 23035
rect 20312 23004 21005 23032
rect 20312 22992 20318 23004
rect 20993 23001 21005 23004
rect 21039 23001 21051 23035
rect 20993 22995 21051 23001
rect 22462 22992 22468 23044
rect 22520 23032 22526 23044
rect 23768 23032 23796 23063
rect 22520 23004 23796 23032
rect 23952 23032 23980 23063
rect 24026 23060 24032 23112
rect 24084 23100 24090 23112
rect 24394 23100 24400 23112
rect 24084 23072 24400 23100
rect 24084 23060 24090 23072
rect 24394 23060 24400 23072
rect 24452 23100 24458 23112
rect 24949 23103 25007 23109
rect 24949 23100 24961 23103
rect 24452 23072 24961 23100
rect 24452 23060 24458 23072
rect 24949 23069 24961 23072
rect 24995 23069 25007 23103
rect 24949 23063 25007 23069
rect 25130 23060 25136 23112
rect 25188 23100 25194 23112
rect 25700 23109 25728 23140
rect 25976 23140 27108 23168
rect 25225 23103 25283 23109
rect 25225 23100 25237 23103
rect 25188 23072 25237 23100
rect 25188 23060 25194 23072
rect 25225 23069 25237 23072
rect 25271 23069 25283 23103
rect 25225 23063 25283 23069
rect 25685 23103 25743 23109
rect 25685 23069 25697 23103
rect 25731 23069 25743 23103
rect 25976 23100 26004 23140
rect 25685 23063 25743 23069
rect 25792 23072 26004 23100
rect 24118 23032 24124 23044
rect 23952 23004 24124 23032
rect 22520 22992 22526 23004
rect 24118 22992 24124 23004
rect 24176 22992 24182 23044
rect 18782 22964 18788 22976
rect 18248 22936 18788 22964
rect 18782 22924 18788 22936
rect 18840 22924 18846 22976
rect 23658 22924 23664 22976
rect 23716 22964 23722 22976
rect 25240 22964 25268 23063
rect 25792 23032 25820 23072
rect 26050 23060 26056 23112
rect 26108 23060 26114 23112
rect 27080 23100 27108 23140
rect 32416 23140 32904 23168
rect 32416 23112 32444 23140
rect 27338 23100 27344 23112
rect 27080 23072 27344 23100
rect 27338 23060 27344 23072
rect 27396 23060 27402 23112
rect 29730 23060 29736 23112
rect 29788 23060 29794 23112
rect 29914 23060 29920 23112
rect 29972 23060 29978 23112
rect 32398 23060 32404 23112
rect 32456 23060 32462 23112
rect 32490 23060 32496 23112
rect 32548 23060 32554 23112
rect 32876 23109 32904 23140
rect 32769 23103 32827 23109
rect 32769 23069 32781 23103
rect 32815 23069 32827 23103
rect 32769 23063 32827 23069
rect 32861 23103 32919 23109
rect 32861 23069 32873 23103
rect 32907 23069 32919 23103
rect 32861 23063 32919 23069
rect 25424 23004 25820 23032
rect 25424 22973 25452 23004
rect 25866 22992 25872 23044
rect 25924 22992 25930 23044
rect 25958 22992 25964 23044
rect 26016 22992 26022 23044
rect 30006 22992 30012 23044
rect 30064 22992 30070 23044
rect 32784 23032 32812 23063
rect 32950 23060 32956 23112
rect 33008 23100 33014 23112
rect 33045 23103 33103 23109
rect 33045 23100 33057 23103
rect 33008 23072 33057 23100
rect 33008 23060 33014 23072
rect 33045 23069 33057 23072
rect 33091 23069 33103 23103
rect 33045 23063 33103 23069
rect 32968 23032 32996 23060
rect 32784 23004 32996 23032
rect 33229 23035 33287 23041
rect 33229 23001 33241 23035
rect 33275 23032 33287 23035
rect 33318 23032 33324 23044
rect 33275 23004 33324 23032
rect 33275 23001 33287 23004
rect 33229 22995 33287 23001
rect 33318 22992 33324 23004
rect 33376 22992 33382 23044
rect 34624 23032 34652 23208
rect 34716 23168 34744 23276
rect 34793 23273 34805 23307
rect 34839 23304 34851 23307
rect 34839 23276 36400 23304
rect 34839 23273 34851 23276
rect 34793 23267 34851 23273
rect 35621 23171 35679 23177
rect 35621 23168 35633 23171
rect 34716 23140 35633 23168
rect 34716 23109 34744 23140
rect 34701 23103 34759 23109
rect 34701 23069 34713 23103
rect 34747 23069 34759 23103
rect 34701 23063 34759 23069
rect 34974 23060 34980 23112
rect 35032 23060 35038 23112
rect 35066 23060 35072 23112
rect 35124 23100 35130 23112
rect 35268 23109 35296 23140
rect 35621 23137 35633 23140
rect 35667 23137 35679 23171
rect 35621 23131 35679 23137
rect 35802 23128 35808 23180
rect 35860 23168 35866 23180
rect 35860 23140 36216 23168
rect 35860 23128 35866 23140
rect 35161 23103 35219 23109
rect 35161 23100 35173 23103
rect 35124 23072 35173 23100
rect 35124 23060 35130 23072
rect 35161 23069 35173 23072
rect 35207 23069 35219 23103
rect 35161 23063 35219 23069
rect 35253 23103 35311 23109
rect 35253 23069 35265 23103
rect 35299 23069 35311 23103
rect 35253 23063 35311 23069
rect 35345 23103 35403 23109
rect 35345 23069 35357 23103
rect 35391 23100 35403 23103
rect 35713 23103 35771 23109
rect 35713 23100 35725 23103
rect 35391 23072 35725 23100
rect 35391 23069 35403 23072
rect 35345 23063 35403 23069
rect 35713 23069 35725 23072
rect 35759 23100 35771 23103
rect 35820 23100 35848 23128
rect 36188 23109 36216 23140
rect 36372 23109 36400 23276
rect 35759 23072 35848 23100
rect 35897 23103 35955 23109
rect 35759 23069 35771 23072
rect 35713 23063 35771 23069
rect 35897 23069 35909 23103
rect 35943 23069 35955 23103
rect 35897 23063 35955 23069
rect 36173 23103 36231 23109
rect 36173 23069 36185 23103
rect 36219 23069 36231 23103
rect 36173 23063 36231 23069
rect 36357 23103 36415 23109
rect 36357 23069 36369 23103
rect 36403 23069 36415 23103
rect 36357 23063 36415 23069
rect 34991 23032 35019 23060
rect 34624 23004 35019 23032
rect 23716 22936 25268 22964
rect 25409 22967 25467 22973
rect 23716 22924 23722 22936
rect 25409 22933 25421 22967
rect 25455 22933 25467 22967
rect 25409 22927 25467 22933
rect 25682 22924 25688 22976
rect 25740 22964 25746 22976
rect 25884 22964 25912 22992
rect 25740 22936 25912 22964
rect 25740 22924 25746 22936
rect 26234 22924 26240 22976
rect 26292 22924 26298 22976
rect 31846 22924 31852 22976
rect 31904 22964 31910 22976
rect 32309 22967 32367 22973
rect 32309 22964 32321 22967
rect 31904 22936 32321 22964
rect 31904 22924 31910 22936
rect 32309 22933 32321 22936
rect 32355 22933 32367 22967
rect 32309 22927 32367 22933
rect 32582 22924 32588 22976
rect 32640 22964 32646 22976
rect 32677 22967 32735 22973
rect 32677 22964 32689 22967
rect 32640 22936 32689 22964
rect 32640 22924 32646 22936
rect 32677 22933 32689 22936
rect 32723 22933 32735 22967
rect 32677 22927 32735 22933
rect 34330 22924 34336 22976
rect 34388 22964 34394 22976
rect 35360 22964 35388 23063
rect 35913 23032 35941 23063
rect 35820 23004 35941 23032
rect 34388 22936 35388 22964
rect 35529 22967 35587 22973
rect 34388 22924 34394 22936
rect 35529 22933 35541 22967
rect 35575 22964 35587 22967
rect 35820 22964 35848 23004
rect 35575 22936 35848 22964
rect 35575 22933 35587 22936
rect 35529 22927 35587 22933
rect 36078 22924 36084 22976
rect 36136 22924 36142 22976
rect 36170 22924 36176 22976
rect 36228 22964 36234 22976
rect 36265 22967 36323 22973
rect 36265 22964 36277 22967
rect 36228 22936 36277 22964
rect 36228 22924 36234 22936
rect 36265 22933 36277 22936
rect 36311 22933 36323 22967
rect 36265 22927 36323 22933
rect 1104 22874 38272 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38272 22874
rect 1104 22800 38272 22822
rect 2682 22720 2688 22772
rect 2740 22760 2746 22772
rect 2869 22763 2927 22769
rect 2869 22760 2881 22763
rect 2740 22732 2881 22760
rect 2740 22720 2746 22732
rect 2869 22729 2881 22732
rect 2915 22729 2927 22763
rect 2869 22723 2927 22729
rect 3142 22720 3148 22772
rect 3200 22760 3206 22772
rect 3421 22763 3479 22769
rect 3421 22760 3433 22763
rect 3200 22732 3433 22760
rect 3200 22720 3206 22732
rect 3421 22729 3433 22732
rect 3467 22729 3479 22763
rect 3421 22723 3479 22729
rect 3970 22720 3976 22772
rect 4028 22720 4034 22772
rect 4430 22720 4436 22772
rect 4488 22760 4494 22772
rect 5077 22763 5135 22769
rect 5077 22760 5089 22763
rect 4488 22732 5089 22760
rect 4488 22720 4494 22732
rect 5077 22729 5089 22732
rect 5123 22729 5135 22763
rect 5537 22763 5595 22769
rect 5537 22760 5549 22763
rect 5077 22723 5135 22729
rect 5184 22732 5549 22760
rect 2498 22652 2504 22704
rect 2556 22692 2562 22704
rect 3050 22692 3056 22704
rect 2556 22664 3056 22692
rect 2556 22652 2562 22664
rect 3050 22652 3056 22664
rect 3108 22692 3114 22704
rect 3605 22695 3663 22701
rect 3605 22692 3617 22695
rect 3108 22664 3617 22692
rect 3108 22652 3114 22664
rect 3605 22661 3617 22664
rect 3651 22692 3663 22695
rect 3651 22664 4108 22692
rect 3651 22661 3663 22664
rect 3605 22655 3663 22661
rect 4080 22636 4108 22664
rect 4522 22652 4528 22704
rect 4580 22692 4586 22704
rect 4798 22692 4804 22704
rect 4580 22664 4804 22692
rect 4580 22652 4586 22664
rect 4798 22652 4804 22664
rect 4856 22692 4862 22704
rect 5184 22692 5212 22732
rect 5537 22729 5549 22732
rect 5583 22729 5595 22763
rect 5537 22723 5595 22729
rect 5626 22720 5632 22772
rect 5684 22720 5690 22772
rect 5828 22732 6684 22760
rect 4856 22664 5212 22692
rect 5445 22695 5503 22701
rect 4856 22652 4862 22664
rect 5445 22661 5457 22695
rect 5491 22692 5503 22695
rect 5644 22692 5672 22720
rect 5491 22664 5672 22692
rect 5491 22661 5503 22664
rect 5445 22655 5503 22661
rect 2777 22627 2835 22633
rect 2777 22593 2789 22627
rect 2823 22593 2835 22627
rect 2777 22587 2835 22593
rect 2792 22556 2820 22587
rect 2958 22584 2964 22636
rect 3016 22584 3022 22636
rect 3789 22627 3847 22633
rect 3789 22593 3801 22627
rect 3835 22624 3847 22627
rect 3878 22624 3884 22636
rect 3835 22596 3884 22624
rect 3835 22593 3847 22596
rect 3789 22587 3847 22593
rect 3878 22584 3884 22596
rect 3936 22584 3942 22636
rect 4062 22584 4068 22636
rect 4120 22584 4126 22636
rect 4706 22584 4712 22636
rect 4764 22624 4770 22636
rect 5166 22624 5172 22636
rect 4764 22596 5172 22624
rect 4764 22584 4770 22596
rect 5166 22584 5172 22596
rect 5224 22624 5230 22636
rect 5261 22627 5319 22633
rect 5261 22624 5273 22627
rect 5224 22596 5273 22624
rect 5224 22584 5230 22596
rect 5261 22593 5273 22596
rect 5307 22624 5319 22627
rect 5537 22627 5595 22633
rect 5537 22624 5549 22627
rect 5307 22596 5549 22624
rect 5307 22593 5319 22596
rect 5261 22587 5319 22593
rect 5537 22593 5549 22596
rect 5583 22593 5595 22627
rect 5644 22624 5672 22664
rect 5721 22627 5779 22633
rect 5721 22624 5733 22627
rect 5644 22596 5733 22624
rect 5537 22587 5595 22593
rect 5721 22593 5733 22596
rect 5767 22593 5779 22627
rect 5721 22587 5779 22593
rect 2866 22556 2872 22568
rect 2792 22528 2872 22556
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 4890 22516 4896 22568
rect 4948 22556 4954 22568
rect 5350 22556 5356 22568
rect 4948 22528 5356 22556
rect 4948 22516 4954 22528
rect 5350 22516 5356 22528
rect 5408 22556 5414 22568
rect 5828 22556 5856 22732
rect 5902 22652 5908 22704
rect 5960 22692 5966 22704
rect 6549 22695 6607 22701
rect 6549 22692 6561 22695
rect 5960 22664 6561 22692
rect 5960 22652 5966 22664
rect 6549 22661 6561 22664
rect 6595 22661 6607 22695
rect 6656 22692 6684 22732
rect 7006 22720 7012 22772
rect 7064 22760 7070 22772
rect 7064 22732 7972 22760
rect 7064 22720 7070 22732
rect 7944 22704 7972 22732
rect 9122 22720 9128 22772
rect 9180 22760 9186 22772
rect 9398 22760 9404 22772
rect 9180 22732 9404 22760
rect 9180 22720 9186 22732
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 9493 22763 9551 22769
rect 9493 22729 9505 22763
rect 9539 22760 9551 22763
rect 9858 22760 9864 22772
rect 9539 22732 9864 22760
rect 9539 22729 9551 22732
rect 9493 22723 9551 22729
rect 9858 22720 9864 22732
rect 9916 22720 9922 22772
rect 11054 22720 11060 22772
rect 11112 22720 11118 22772
rect 11517 22763 11575 22769
rect 11517 22729 11529 22763
rect 11563 22729 11575 22763
rect 11517 22723 11575 22729
rect 11885 22763 11943 22769
rect 11885 22729 11897 22763
rect 11931 22760 11943 22763
rect 12342 22760 12348 22772
rect 11931 22732 12348 22760
rect 11931 22729 11943 22732
rect 11885 22723 11943 22729
rect 7374 22692 7380 22704
rect 6656 22664 7380 22692
rect 6549 22655 6607 22661
rect 7374 22652 7380 22664
rect 7432 22652 7438 22704
rect 7650 22652 7656 22704
rect 7708 22652 7714 22704
rect 7926 22652 7932 22704
rect 7984 22692 7990 22704
rect 8021 22695 8079 22701
rect 8021 22692 8033 22695
rect 7984 22664 8033 22692
rect 7984 22652 7990 22664
rect 8021 22661 8033 22664
rect 8067 22661 8079 22695
rect 8021 22655 8079 22661
rect 8205 22695 8263 22701
rect 8205 22661 8217 22695
rect 8251 22692 8263 22695
rect 11330 22692 11336 22704
rect 8251 22664 11336 22692
rect 8251 22661 8263 22664
rect 8205 22655 8263 22661
rect 11330 22652 11336 22664
rect 11388 22652 11394 22704
rect 6365 22627 6423 22633
rect 6365 22593 6377 22627
rect 6411 22624 6423 22627
rect 6914 22624 6920 22636
rect 6411 22596 6920 22624
rect 6411 22593 6423 22596
rect 6365 22587 6423 22593
rect 6914 22584 6920 22596
rect 6972 22584 6978 22636
rect 5408 22528 5856 22556
rect 6733 22559 6791 22565
rect 5408 22516 5414 22528
rect 6733 22525 6745 22559
rect 6779 22556 6791 22559
rect 7668 22556 7696 22652
rect 7837 22627 7895 22633
rect 7837 22593 7849 22627
rect 7883 22624 7895 22627
rect 8110 22624 8116 22636
rect 7883 22596 8116 22624
rect 7883 22593 7895 22596
rect 7837 22587 7895 22593
rect 8110 22584 8116 22596
rect 8168 22584 8174 22636
rect 8754 22584 8760 22636
rect 8812 22624 8818 22636
rect 9677 22627 9735 22633
rect 9677 22624 9689 22627
rect 8812 22596 9689 22624
rect 8812 22584 8818 22596
rect 9677 22593 9689 22596
rect 9723 22624 9735 22627
rect 9861 22627 9919 22633
rect 9723 22596 9812 22624
rect 9723 22593 9735 22596
rect 9677 22587 9735 22593
rect 6779 22528 7696 22556
rect 6779 22525 6791 22528
rect 6733 22519 6791 22525
rect 3602 22448 3608 22500
rect 3660 22488 3666 22500
rect 6270 22488 6276 22500
rect 3660 22460 6276 22488
rect 3660 22448 3666 22460
rect 6270 22448 6276 22460
rect 6328 22448 6334 22500
rect 9784 22488 9812 22596
rect 9861 22593 9873 22627
rect 9907 22624 9919 22627
rect 10134 22624 10140 22636
rect 9907 22596 10140 22624
rect 9907 22593 9919 22596
rect 9861 22587 9919 22593
rect 10134 22584 10140 22596
rect 10192 22584 10198 22636
rect 11241 22627 11299 22633
rect 11241 22593 11253 22627
rect 11287 22624 11299 22627
rect 11532 22624 11560 22723
rect 12342 22720 12348 22732
rect 12400 22720 12406 22772
rect 12434 22720 12440 22772
rect 12492 22760 12498 22772
rect 12989 22763 13047 22769
rect 12989 22760 13001 22763
rect 12492 22732 13001 22760
rect 12492 22720 12498 22732
rect 12989 22729 13001 22732
rect 13035 22729 13047 22763
rect 12989 22723 13047 22729
rect 13817 22763 13875 22769
rect 13817 22729 13829 22763
rect 13863 22760 13875 22763
rect 14090 22760 14096 22772
rect 13863 22732 14096 22760
rect 13863 22729 13875 22732
rect 13817 22723 13875 22729
rect 14090 22720 14096 22732
rect 14148 22720 14154 22772
rect 15194 22720 15200 22772
rect 15252 22760 15258 22772
rect 15289 22763 15347 22769
rect 15289 22760 15301 22763
rect 15252 22732 15301 22760
rect 15252 22720 15258 22732
rect 15289 22729 15301 22732
rect 15335 22729 15347 22763
rect 15289 22723 15347 22729
rect 15470 22720 15476 22772
rect 15528 22720 15534 22772
rect 15838 22720 15844 22772
rect 15896 22760 15902 22772
rect 17957 22763 18015 22769
rect 15896 22732 16160 22760
rect 15896 22720 15902 22732
rect 16132 22704 16160 22732
rect 17957 22729 17969 22763
rect 18003 22760 18015 22763
rect 18506 22760 18512 22772
rect 18003 22732 18512 22760
rect 18003 22729 18015 22732
rect 17957 22723 18015 22729
rect 18506 22720 18512 22732
rect 18564 22720 18570 22772
rect 20438 22720 20444 22772
rect 20496 22720 20502 22772
rect 22097 22763 22155 22769
rect 22097 22729 22109 22763
rect 22143 22760 22155 22763
rect 22922 22760 22928 22772
rect 22143 22732 22928 22760
rect 22143 22729 22155 22732
rect 22097 22723 22155 22729
rect 22922 22720 22928 22732
rect 22980 22720 22986 22772
rect 23658 22760 23664 22772
rect 23032 22732 23664 22760
rect 13633 22695 13691 22701
rect 13633 22661 13645 22695
rect 13679 22692 13691 22695
rect 13998 22692 14004 22704
rect 13679 22664 14004 22692
rect 13679 22661 13691 22664
rect 13633 22655 13691 22661
rect 13998 22652 14004 22664
rect 14056 22692 14062 22704
rect 14056 22664 14320 22692
rect 14056 22652 14062 22664
rect 11287 22596 11560 22624
rect 12345 22627 12403 22633
rect 11287 22593 11299 22596
rect 11241 22587 11299 22593
rect 12345 22593 12357 22627
rect 12391 22624 12403 22627
rect 12434 22624 12440 22636
rect 12391 22596 12440 22624
rect 12391 22593 12403 22596
rect 12345 22587 12403 22593
rect 9953 22559 10011 22565
rect 9953 22525 9965 22559
rect 9999 22556 10011 22559
rect 10042 22556 10048 22568
rect 9999 22528 10048 22556
rect 9999 22525 10011 22528
rect 9953 22519 10011 22525
rect 10042 22516 10048 22528
rect 10100 22516 10106 22568
rect 11974 22516 11980 22568
rect 12032 22516 12038 22568
rect 12158 22516 12164 22568
rect 12216 22516 12222 22568
rect 12176 22488 12204 22516
rect 9784 22460 12204 22488
rect 3694 22380 3700 22432
rect 3752 22420 3758 22432
rect 4154 22420 4160 22432
rect 3752 22392 4160 22420
rect 3752 22380 3758 22392
rect 4154 22380 4160 22392
rect 4212 22420 4218 22432
rect 6178 22420 6184 22432
rect 4212 22392 6184 22420
rect 4212 22380 4218 22392
rect 6178 22380 6184 22392
rect 6236 22420 6242 22432
rect 12360 22420 12388 22587
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 12526 22584 12532 22636
rect 12584 22584 12590 22636
rect 12621 22627 12679 22633
rect 12621 22593 12633 22627
rect 12667 22593 12679 22627
rect 12621 22587 12679 22593
rect 12713 22627 12771 22633
rect 12713 22593 12725 22627
rect 12759 22624 12771 22627
rect 13357 22627 13415 22633
rect 12759 22596 13308 22624
rect 12759 22593 12771 22596
rect 12713 22587 12771 22593
rect 12636 22556 12664 22587
rect 12802 22556 12808 22568
rect 12636 22528 12808 22556
rect 12802 22516 12808 22528
rect 12860 22516 12866 22568
rect 13280 22488 13308 22596
rect 13357 22593 13369 22627
rect 13403 22624 13415 22627
rect 13446 22624 13452 22636
rect 13403 22596 13452 22624
rect 13403 22593 13415 22596
rect 13357 22587 13415 22593
rect 13446 22584 13452 22596
rect 13504 22584 13510 22636
rect 13541 22627 13599 22633
rect 13541 22593 13553 22627
rect 13587 22624 13599 22627
rect 14182 22624 14188 22636
rect 13587 22596 14188 22624
rect 13587 22593 13599 22596
rect 13541 22587 13599 22593
rect 14182 22584 14188 22596
rect 14240 22584 14246 22636
rect 14292 22633 14320 22664
rect 16114 22652 16120 22704
rect 16172 22652 16178 22704
rect 16301 22695 16359 22701
rect 16301 22661 16313 22695
rect 16347 22692 16359 22695
rect 16758 22692 16764 22704
rect 16347 22664 16764 22692
rect 16347 22661 16359 22664
rect 16301 22655 16359 22661
rect 16758 22652 16764 22664
rect 16816 22652 16822 22704
rect 17494 22652 17500 22704
rect 17552 22692 17558 22704
rect 19334 22692 19340 22704
rect 17552 22664 19340 22692
rect 17552 22652 17558 22664
rect 19334 22652 19340 22664
rect 19392 22652 19398 22704
rect 23032 22692 23060 22732
rect 23658 22720 23664 22732
rect 23716 22720 23722 22772
rect 23750 22720 23756 22772
rect 23808 22760 23814 22772
rect 24397 22763 24455 22769
rect 24397 22760 24409 22763
rect 23808 22732 24409 22760
rect 23808 22720 23814 22732
rect 24397 22729 24409 22732
rect 24443 22729 24455 22763
rect 24397 22723 24455 22729
rect 25590 22720 25596 22772
rect 25648 22720 25654 22772
rect 26234 22720 26240 22772
rect 26292 22720 26298 22772
rect 27522 22720 27528 22772
rect 27580 22720 27586 22772
rect 27985 22763 28043 22769
rect 27985 22729 27997 22763
rect 28031 22760 28043 22763
rect 28350 22760 28356 22772
rect 28031 22732 28356 22760
rect 28031 22729 28043 22732
rect 27985 22723 28043 22729
rect 28350 22720 28356 22732
rect 28408 22720 28414 22772
rect 29914 22720 29920 22772
rect 29972 22760 29978 22772
rect 30285 22763 30343 22769
rect 30285 22760 30297 22763
rect 29972 22732 30297 22760
rect 29972 22720 29978 22732
rect 30285 22729 30297 22732
rect 30331 22729 30343 22763
rect 30285 22723 30343 22729
rect 32217 22763 32275 22769
rect 32217 22729 32229 22763
rect 32263 22760 32275 22763
rect 32490 22760 32496 22772
rect 32263 22732 32496 22760
rect 32263 22729 32275 22732
rect 32217 22723 32275 22729
rect 32490 22720 32496 22732
rect 32548 22720 32554 22772
rect 33042 22720 33048 22772
rect 33100 22760 33106 22772
rect 33689 22763 33747 22769
rect 33689 22760 33701 22763
rect 33100 22732 33701 22760
rect 33100 22720 33106 22732
rect 33689 22729 33701 22732
rect 33735 22729 33747 22763
rect 33689 22723 33747 22729
rect 35066 22720 35072 22772
rect 35124 22760 35130 22772
rect 35124 22732 36400 22760
rect 35124 22720 35130 22732
rect 25608 22692 25636 22720
rect 26252 22692 26280 22720
rect 35161 22695 35219 22701
rect 22020 22664 22600 22692
rect 14277 22627 14335 22633
rect 14277 22593 14289 22627
rect 14323 22593 14335 22627
rect 14277 22587 14335 22593
rect 14458 22584 14464 22636
rect 14516 22624 14522 22636
rect 14642 22624 14648 22636
rect 14516 22596 14648 22624
rect 14516 22584 14522 22596
rect 14642 22584 14648 22596
rect 14700 22584 14706 22636
rect 15471 22627 15529 22633
rect 15471 22593 15483 22627
rect 15517 22624 15529 22627
rect 15562 22624 15568 22636
rect 15517 22596 15568 22624
rect 15517 22593 15529 22596
rect 15471 22587 15529 22593
rect 15562 22584 15568 22596
rect 15620 22584 15626 22636
rect 15933 22627 15991 22633
rect 15933 22593 15945 22627
rect 15979 22624 15991 22627
rect 15979 22596 16344 22624
rect 15979 22593 15991 22596
rect 15933 22587 15991 22593
rect 16316 22568 16344 22596
rect 16850 22584 16856 22636
rect 16908 22624 16914 22636
rect 17126 22624 17132 22636
rect 16908 22596 17132 22624
rect 16908 22584 16914 22596
rect 17126 22584 17132 22596
rect 17184 22584 17190 22636
rect 17310 22584 17316 22636
rect 17368 22584 17374 22636
rect 17862 22584 17868 22636
rect 17920 22584 17926 22636
rect 20714 22584 20720 22636
rect 20772 22584 20778 22636
rect 21910 22584 21916 22636
rect 21968 22624 21974 22636
rect 22020 22633 22048 22664
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21968 22596 22017 22624
rect 21968 22584 21974 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 22186 22584 22192 22636
rect 22244 22624 22250 22636
rect 22462 22624 22468 22636
rect 22244 22596 22468 22624
rect 22244 22584 22250 22596
rect 22462 22584 22468 22596
rect 22520 22584 22526 22636
rect 22572 22633 22600 22664
rect 22664 22664 23060 22692
rect 23308 22664 24532 22692
rect 22664 22633 22692 22664
rect 23308 22636 23336 22664
rect 22557 22627 22615 22633
rect 22557 22593 22569 22627
rect 22603 22593 22615 22627
rect 22557 22587 22615 22593
rect 22649 22627 22707 22633
rect 22649 22593 22661 22627
rect 22695 22593 22707 22627
rect 22649 22587 22707 22593
rect 23017 22627 23075 22633
rect 23017 22593 23029 22627
rect 23063 22624 23075 22627
rect 23290 22624 23296 22636
rect 23063 22596 23296 22624
rect 23063 22593 23075 22596
rect 23017 22587 23075 22593
rect 14660 22528 15976 22556
rect 14660 22488 14688 22528
rect 15841 22491 15899 22497
rect 15841 22488 15853 22491
rect 13280 22460 14688 22488
rect 15120 22460 15853 22488
rect 6236 22392 12388 22420
rect 6236 22380 6242 22392
rect 14182 22380 14188 22432
rect 14240 22420 14246 22432
rect 15120 22420 15148 22460
rect 15841 22457 15853 22460
rect 15887 22457 15899 22491
rect 15841 22451 15899 22457
rect 14240 22392 15148 22420
rect 15948 22420 15976 22528
rect 16298 22516 16304 22568
rect 16356 22516 16362 22568
rect 16485 22559 16543 22565
rect 16485 22525 16497 22559
rect 16531 22556 16543 22559
rect 17328 22556 17356 22584
rect 16531 22528 17356 22556
rect 16531 22525 16543 22528
rect 16485 22519 16543 22525
rect 17494 22516 17500 22568
rect 17552 22556 17558 22568
rect 22572 22556 22600 22587
rect 23290 22584 23296 22596
rect 23348 22584 23354 22636
rect 23382 22584 23388 22636
rect 23440 22584 23446 22636
rect 23566 22584 23572 22636
rect 23624 22584 23630 22636
rect 24026 22584 24032 22636
rect 24084 22584 24090 22636
rect 24504 22633 24532 22664
rect 25608 22664 26193 22692
rect 26252 22664 30696 22692
rect 25608 22633 25636 22664
rect 26165 22636 26193 22664
rect 24305 22627 24363 22633
rect 24305 22593 24317 22627
rect 24351 22593 24363 22627
rect 24305 22587 24363 22593
rect 24489 22627 24547 22633
rect 24489 22593 24501 22627
rect 24535 22593 24547 22627
rect 24489 22587 24547 22593
rect 25593 22627 25651 22633
rect 25593 22593 25605 22627
rect 25639 22593 25651 22627
rect 25593 22587 25651 22593
rect 24118 22556 24124 22568
rect 17552 22528 22508 22556
rect 22572 22528 24124 22556
rect 17552 22516 17558 22528
rect 16022 22448 16028 22500
rect 16080 22488 16086 22500
rect 16758 22488 16764 22500
rect 16080 22460 16764 22488
rect 16080 22448 16086 22460
rect 16758 22448 16764 22460
rect 16816 22448 16822 22500
rect 19242 22448 19248 22500
rect 19300 22488 19306 22500
rect 20070 22488 20076 22500
rect 19300 22460 20076 22488
rect 19300 22448 19306 22460
rect 20070 22448 20076 22460
rect 20128 22448 20134 22500
rect 21818 22420 21824 22432
rect 15948 22392 21824 22420
rect 14240 22380 14246 22392
rect 21818 22380 21824 22392
rect 21876 22380 21882 22432
rect 22480 22420 22508 22528
rect 24118 22516 24124 22528
rect 24176 22556 24182 22568
rect 24320 22556 24348 22587
rect 25774 22584 25780 22636
rect 25832 22584 25838 22636
rect 26142 22584 26148 22636
rect 26200 22624 26206 22636
rect 26510 22624 26516 22636
rect 26200 22596 26516 22624
rect 26200 22584 26206 22596
rect 26510 22584 26516 22596
rect 26568 22584 26574 22636
rect 26602 22584 26608 22636
rect 26660 22624 26666 22636
rect 26973 22627 27031 22633
rect 26973 22624 26985 22627
rect 26660 22596 26985 22624
rect 26660 22584 26666 22596
rect 26973 22593 26985 22596
rect 27019 22593 27031 22627
rect 26973 22587 27031 22593
rect 27154 22584 27160 22636
rect 27212 22584 27218 22636
rect 27249 22627 27307 22633
rect 27249 22593 27261 22627
rect 27295 22593 27307 22627
rect 27249 22587 27307 22593
rect 27341 22627 27399 22633
rect 27341 22593 27353 22627
rect 27387 22624 27399 22627
rect 27430 22624 27436 22636
rect 27387 22596 27436 22624
rect 27387 22593 27399 22596
rect 27341 22587 27399 22593
rect 24176 22528 24348 22556
rect 24176 22516 24182 22528
rect 25866 22516 25872 22568
rect 25924 22556 25930 22568
rect 27264 22556 27292 22587
rect 25924 22528 27292 22556
rect 25924 22516 25930 22528
rect 23934 22448 23940 22500
rect 23992 22448 23998 22500
rect 26050 22448 26056 22500
rect 26108 22488 26114 22500
rect 27356 22488 27384 22587
rect 27430 22584 27436 22596
rect 27488 22584 27494 22636
rect 27706 22584 27712 22636
rect 27764 22584 27770 22636
rect 29656 22633 29684 22664
rect 29641 22627 29699 22633
rect 29641 22593 29653 22627
rect 29687 22593 29699 22627
rect 29641 22587 29699 22593
rect 29825 22627 29883 22633
rect 29825 22593 29837 22627
rect 29871 22624 29883 22627
rect 29917 22627 29975 22633
rect 29917 22624 29929 22627
rect 29871 22596 29929 22624
rect 29871 22593 29883 22596
rect 29825 22587 29883 22593
rect 29917 22593 29929 22596
rect 29963 22624 29975 22627
rect 30190 22624 30196 22636
rect 29963 22596 30196 22624
rect 29963 22593 29975 22596
rect 29917 22587 29975 22593
rect 30190 22584 30196 22596
rect 30248 22584 30254 22636
rect 30392 22633 30420 22664
rect 30668 22633 30696 22664
rect 32140 22664 33180 22692
rect 32140 22636 32168 22664
rect 30377 22627 30435 22633
rect 30377 22593 30389 22627
rect 30423 22593 30435 22627
rect 30377 22587 30435 22593
rect 30469 22627 30527 22633
rect 30469 22593 30481 22627
rect 30515 22593 30527 22627
rect 30469 22587 30527 22593
rect 30653 22627 30711 22633
rect 30653 22593 30665 22627
rect 30699 22593 30711 22627
rect 30653 22587 30711 22593
rect 30009 22559 30067 22565
rect 30009 22525 30021 22559
rect 30055 22556 30067 22559
rect 30484 22556 30512 22587
rect 32122 22584 32128 22636
rect 32180 22584 32186 22636
rect 32309 22627 32367 22633
rect 32309 22593 32321 22627
rect 32355 22624 32367 22627
rect 32398 22624 32404 22636
rect 32355 22596 32404 22624
rect 32355 22593 32367 22596
rect 32309 22587 32367 22593
rect 32398 22584 32404 22596
rect 32456 22584 32462 22636
rect 32770 22627 32828 22633
rect 32770 22593 32782 22627
rect 32816 22622 32828 22627
rect 33042 22624 33048 22636
rect 32876 22622 33048 22624
rect 32816 22596 33048 22622
rect 32816 22594 32904 22596
rect 32816 22593 32828 22594
rect 32770 22587 32828 22593
rect 33042 22584 33048 22596
rect 33100 22584 33106 22636
rect 33152 22633 33180 22664
rect 35161 22661 35173 22695
rect 35207 22692 35219 22695
rect 36170 22692 36176 22704
rect 35207 22664 36176 22692
rect 35207 22661 35219 22664
rect 35161 22655 35219 22661
rect 36170 22652 36176 22664
rect 36228 22652 36234 22704
rect 36372 22692 36400 22732
rect 36446 22720 36452 22772
rect 36504 22760 36510 22772
rect 37369 22763 37427 22769
rect 37369 22760 37381 22763
rect 36504 22732 37381 22760
rect 36504 22720 36510 22732
rect 37369 22729 37381 22732
rect 37415 22729 37427 22763
rect 37369 22723 37427 22729
rect 36817 22695 36875 22701
rect 36817 22692 36829 22695
rect 36372 22664 36829 22692
rect 33137 22627 33195 22633
rect 33137 22593 33149 22627
rect 33183 22593 33195 22627
rect 33137 22587 33195 22593
rect 33226 22584 33232 22636
rect 33284 22584 33290 22636
rect 33318 22584 33324 22636
rect 33376 22624 33382 22636
rect 33413 22627 33471 22633
rect 33413 22624 33425 22627
rect 33376 22596 33425 22624
rect 33376 22584 33382 22596
rect 33413 22593 33425 22596
rect 33459 22593 33471 22627
rect 33413 22587 33471 22593
rect 33505 22627 33563 22633
rect 33505 22593 33517 22627
rect 33551 22624 33563 22627
rect 34422 22624 34428 22636
rect 33551 22596 34428 22624
rect 33551 22593 33563 22596
rect 33505 22587 33563 22593
rect 34422 22584 34428 22596
rect 34480 22584 34486 22636
rect 34974 22584 34980 22636
rect 35032 22584 35038 22636
rect 35342 22584 35348 22636
rect 35400 22584 35406 22636
rect 35437 22627 35495 22633
rect 35437 22593 35449 22627
rect 35483 22624 35495 22627
rect 35802 22624 35808 22636
rect 35483 22596 35808 22624
rect 35483 22593 35495 22596
rect 35437 22587 35495 22593
rect 35802 22584 35808 22596
rect 35860 22584 35866 22636
rect 36081 22627 36139 22633
rect 36081 22593 36093 22627
rect 36127 22593 36139 22627
rect 36081 22587 36139 22593
rect 30055 22528 30512 22556
rect 30055 22525 30067 22528
rect 30009 22519 30067 22525
rect 31846 22516 31852 22568
rect 31904 22556 31910 22568
rect 32677 22559 32735 22565
rect 32677 22556 32689 22559
rect 31904 22528 32689 22556
rect 31904 22516 31910 22528
rect 32677 22525 32689 22528
rect 32723 22525 32735 22559
rect 32677 22519 32735 22525
rect 32861 22559 32919 22565
rect 32861 22525 32873 22559
rect 32907 22525 32919 22559
rect 32861 22519 32919 22525
rect 26108 22460 27384 22488
rect 32876 22488 32904 22519
rect 32950 22516 32956 22568
rect 33008 22516 33014 22568
rect 34992 22556 35020 22584
rect 36096 22556 36124 22587
rect 36262 22584 36268 22636
rect 36320 22584 36326 22636
rect 36372 22633 36400 22664
rect 36817 22661 36829 22664
rect 36863 22692 36875 22695
rect 36863 22664 37320 22692
rect 36863 22661 36875 22664
rect 36817 22655 36875 22661
rect 37292 22633 37320 22664
rect 36357 22627 36415 22633
rect 36357 22593 36369 22627
rect 36403 22593 36415 22627
rect 36541 22627 36599 22633
rect 36541 22624 36553 22627
rect 36357 22587 36415 22593
rect 36464 22596 36553 22624
rect 34992 22528 36124 22556
rect 33226 22488 33232 22500
rect 32876 22460 33232 22488
rect 26108 22448 26114 22460
rect 33226 22448 33232 22460
rect 33284 22448 33290 22500
rect 36096 22488 36124 22528
rect 36464 22488 36492 22596
rect 36541 22593 36553 22596
rect 36587 22624 36599 22627
rect 36633 22627 36691 22633
rect 36633 22624 36645 22627
rect 36587 22596 36645 22624
rect 36587 22593 36599 22596
rect 36541 22587 36599 22593
rect 36633 22593 36645 22596
rect 36679 22593 36691 22627
rect 36633 22587 36691 22593
rect 37277 22627 37335 22633
rect 37277 22593 37289 22627
rect 37323 22593 37335 22627
rect 37277 22587 37335 22593
rect 37550 22584 37556 22636
rect 37608 22624 37614 22636
rect 37645 22627 37703 22633
rect 37645 22624 37657 22627
rect 37608 22596 37657 22624
rect 37608 22584 37614 22596
rect 37645 22593 37657 22596
rect 37691 22593 37703 22627
rect 37645 22587 37703 22593
rect 36096 22460 36492 22488
rect 37826 22448 37832 22500
rect 37884 22448 37890 22500
rect 24762 22420 24768 22432
rect 22480 22392 24768 22420
rect 24762 22380 24768 22392
rect 24820 22380 24826 22432
rect 25409 22423 25467 22429
rect 25409 22389 25421 22423
rect 25455 22420 25467 22423
rect 25958 22420 25964 22432
rect 25455 22392 25964 22420
rect 25455 22389 25467 22392
rect 25409 22383 25467 22389
rect 25958 22380 25964 22392
rect 26016 22380 26022 22432
rect 29457 22423 29515 22429
rect 29457 22389 29469 22423
rect 29503 22420 29515 22423
rect 29730 22420 29736 22432
rect 29503 22392 29736 22420
rect 29503 22389 29515 22392
rect 29457 22383 29515 22389
rect 29730 22380 29736 22392
rect 29788 22380 29794 22432
rect 30650 22380 30656 22432
rect 30708 22380 30714 22432
rect 32490 22380 32496 22432
rect 32548 22380 32554 22432
rect 32582 22380 32588 22432
rect 32640 22420 32646 22432
rect 34790 22420 34796 22432
rect 32640 22392 34796 22420
rect 32640 22380 32646 22392
rect 34790 22380 34796 22392
rect 34848 22420 34854 22432
rect 35161 22423 35219 22429
rect 35161 22420 35173 22423
rect 34848 22392 35173 22420
rect 34848 22380 34854 22392
rect 35161 22389 35173 22392
rect 35207 22389 35219 22423
rect 35161 22383 35219 22389
rect 35894 22380 35900 22432
rect 35952 22420 35958 22432
rect 36081 22423 36139 22429
rect 36081 22420 36093 22423
rect 35952 22392 36093 22420
rect 35952 22380 35958 22392
rect 36081 22389 36093 22392
rect 36127 22389 36139 22423
rect 36081 22383 36139 22389
rect 36446 22380 36452 22432
rect 36504 22380 36510 22432
rect 36998 22380 37004 22432
rect 37056 22380 37062 22432
rect 1104 22330 38272 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38272 22330
rect 1104 22256 38272 22278
rect 3602 22176 3608 22228
rect 3660 22216 3666 22228
rect 3973 22219 4031 22225
rect 3973 22216 3985 22219
rect 3660 22188 3985 22216
rect 3660 22176 3666 22188
rect 3973 22185 3985 22188
rect 4019 22185 4031 22219
rect 3973 22179 4031 22185
rect 9674 22176 9680 22228
rect 9732 22216 9738 22228
rect 10321 22219 10379 22225
rect 10321 22216 10333 22219
rect 9732 22188 10333 22216
rect 9732 22176 9738 22188
rect 10321 22185 10333 22188
rect 10367 22185 10379 22219
rect 10321 22179 10379 22185
rect 11974 22176 11980 22228
rect 12032 22216 12038 22228
rect 12161 22219 12219 22225
rect 12161 22216 12173 22219
rect 12032 22188 12173 22216
rect 12032 22176 12038 22188
rect 12161 22185 12173 22188
rect 12207 22185 12219 22219
rect 25866 22216 25872 22228
rect 12161 22179 12219 22185
rect 12406 22188 25872 22216
rect 4157 22151 4215 22157
rect 4157 22117 4169 22151
rect 4203 22148 4215 22151
rect 5994 22148 6000 22160
rect 4203 22120 6000 22148
rect 4203 22117 4215 22120
rect 4157 22111 4215 22117
rect 1946 21972 1952 22024
rect 2004 21972 2010 22024
rect 4062 22012 4068 22024
rect 3804 21984 4068 22012
rect 3804 21953 3832 21984
rect 4062 21972 4068 21984
rect 4120 21972 4126 22024
rect 4172 22012 4200 22111
rect 5994 22108 6000 22120
rect 6052 22108 6058 22160
rect 6270 22108 6276 22160
rect 6328 22148 6334 22160
rect 12406 22148 12434 22188
rect 25866 22176 25872 22188
rect 25924 22176 25930 22228
rect 27356 22188 28212 22216
rect 6328 22120 12434 22148
rect 6328 22108 6334 22120
rect 15378 22108 15384 22160
rect 15436 22148 15442 22160
rect 16390 22148 16396 22160
rect 15436 22120 16396 22148
rect 15436 22108 15442 22120
rect 16390 22108 16396 22120
rect 16448 22108 16454 22160
rect 16758 22108 16764 22160
rect 16816 22148 16822 22160
rect 16816 22120 16896 22148
rect 16816 22108 16822 22120
rect 10042 22040 10048 22092
rect 10100 22040 10106 22092
rect 11609 22083 11667 22089
rect 11609 22049 11621 22083
rect 11655 22049 11667 22083
rect 11609 22043 11667 22049
rect 4249 22015 4307 22021
rect 4249 22012 4261 22015
rect 4172 21984 4261 22012
rect 4249 21981 4261 21984
rect 4295 21981 4307 22015
rect 4249 21975 4307 21981
rect 7745 22015 7803 22021
rect 7745 21981 7757 22015
rect 7791 21981 7803 22015
rect 10060 22012 10088 22040
rect 10229 22015 10287 22021
rect 10229 22012 10241 22015
rect 10060 21984 10241 22012
rect 7745 21975 7803 21981
rect 10229 21981 10241 21984
rect 10275 21981 10287 22015
rect 10229 21975 10287 21981
rect 10413 22015 10471 22021
rect 10413 21981 10425 22015
rect 10459 22012 10471 22015
rect 11422 22012 11428 22024
rect 10459 21984 11428 22012
rect 10459 21981 10471 21984
rect 10413 21975 10471 21981
rect 3789 21947 3847 21953
rect 3789 21913 3801 21947
rect 3835 21913 3847 21947
rect 3789 21907 3847 21913
rect 3878 21904 3884 21956
rect 3936 21904 3942 21956
rect 7760 21944 7788 21975
rect 5828 21916 7788 21944
rect 10244 21944 10272 21975
rect 11422 21972 11428 21984
rect 11480 21972 11486 22024
rect 11624 21944 11652 22043
rect 12158 22040 12164 22092
rect 12216 22080 12222 22092
rect 12253 22083 12311 22089
rect 12253 22080 12265 22083
rect 12216 22052 12265 22080
rect 12216 22040 12222 22052
rect 12253 22049 12265 22052
rect 12299 22049 12311 22083
rect 12253 22043 12311 22049
rect 14366 22040 14372 22092
rect 14424 22080 14430 22092
rect 14461 22083 14519 22089
rect 14461 22080 14473 22083
rect 14424 22052 14473 22080
rect 14424 22040 14430 22052
rect 14461 22049 14473 22052
rect 14507 22049 14519 22083
rect 15654 22080 15660 22092
rect 14461 22043 14519 22049
rect 15396 22052 15660 22080
rect 15396 22024 15424 22052
rect 15654 22040 15660 22052
rect 15712 22080 15718 22092
rect 16485 22083 16543 22089
rect 16485 22080 16497 22083
rect 15712 22052 15884 22080
rect 15712 22040 15718 22052
rect 12805 22015 12863 22021
rect 12805 21981 12817 22015
rect 12851 22012 12863 22015
rect 13722 22012 13728 22024
rect 12851 21984 13728 22012
rect 12851 21981 12863 21984
rect 12805 21975 12863 21981
rect 13722 21972 13728 21984
rect 13780 21972 13786 22024
rect 14182 21972 14188 22024
rect 14240 22012 14246 22024
rect 14829 22015 14887 22021
rect 14829 22012 14841 22015
rect 14240 21984 14841 22012
rect 14240 21972 14246 21984
rect 14829 21981 14841 21984
rect 14875 21981 14887 22015
rect 14829 21975 14887 21981
rect 15013 22015 15071 22021
rect 15013 21981 15025 22015
rect 15059 21981 15071 22015
rect 15013 21975 15071 21981
rect 12437 21947 12495 21953
rect 10244 21916 12204 21944
rect 1762 21836 1768 21888
rect 1820 21836 1826 21888
rect 3896 21876 3924 21904
rect 5828 21888 5856 21916
rect 12176 21888 12204 21916
rect 12437 21913 12449 21947
rect 12483 21944 12495 21947
rect 14550 21944 14556 21956
rect 12483 21916 14556 21944
rect 12483 21913 12495 21916
rect 12437 21907 12495 21913
rect 14550 21904 14556 21916
rect 14608 21904 14614 21956
rect 15028 21944 15056 21975
rect 15378 21972 15384 22024
rect 15436 21972 15442 22024
rect 15470 21972 15476 22024
rect 15528 21972 15534 22024
rect 15562 21972 15568 22024
rect 15620 21972 15626 22024
rect 15856 22021 15884 22052
rect 16316 22052 16497 22080
rect 16316 22024 16344 22052
rect 16485 22049 16497 22052
rect 16531 22049 16543 22083
rect 16868 22080 16896 22120
rect 16942 22108 16948 22160
rect 17000 22148 17006 22160
rect 17037 22151 17095 22157
rect 17037 22148 17049 22151
rect 17000 22120 17049 22148
rect 17000 22108 17006 22120
rect 17037 22117 17049 22120
rect 17083 22117 17095 22151
rect 17037 22111 17095 22117
rect 17218 22108 17224 22160
rect 17276 22148 17282 22160
rect 17862 22148 17868 22160
rect 17276 22120 17868 22148
rect 17276 22108 17282 22120
rect 17862 22108 17868 22120
rect 17920 22108 17926 22160
rect 19242 22108 19248 22160
rect 19300 22108 19306 22160
rect 23566 22108 23572 22160
rect 23624 22148 23630 22160
rect 24213 22151 24271 22157
rect 24213 22148 24225 22151
rect 23624 22120 24225 22148
rect 23624 22108 23630 22120
rect 24213 22117 24225 22120
rect 24259 22148 24271 22151
rect 24578 22148 24584 22160
rect 24259 22120 24584 22148
rect 24259 22117 24271 22120
rect 24213 22111 24271 22117
rect 24578 22108 24584 22120
rect 24636 22108 24642 22160
rect 24946 22108 24952 22160
rect 25004 22148 25010 22160
rect 27356 22148 27384 22188
rect 27801 22151 27859 22157
rect 27801 22148 27813 22151
rect 25004 22120 27384 22148
rect 27448 22120 27813 22148
rect 25004 22108 25010 22120
rect 23661 22083 23719 22089
rect 16868 22052 19840 22080
rect 16485 22043 16543 22049
rect 15841 22015 15899 22021
rect 15841 21981 15853 22015
rect 15887 21981 15899 22015
rect 15841 21975 15899 21981
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 22012 16083 22015
rect 16114 22012 16120 22024
rect 16071 21984 16120 22012
rect 16071 21981 16083 21984
rect 16025 21975 16083 21981
rect 16114 21972 16120 21984
rect 16172 21972 16178 22024
rect 16298 21972 16304 22024
rect 16356 21972 16362 22024
rect 16390 21972 16396 22024
rect 16448 22012 16454 22024
rect 16758 22012 16764 22024
rect 16448 21984 16764 22012
rect 16448 21972 16454 21984
rect 16758 21972 16764 21984
rect 16816 21972 16822 22024
rect 16853 22015 16911 22021
rect 16853 21981 16865 22015
rect 16899 21981 16911 22015
rect 16853 21975 16911 21981
rect 15102 21944 15108 21956
rect 15028 21916 15108 21944
rect 15102 21904 15108 21916
rect 15160 21944 15166 21956
rect 16316 21944 16344 21972
rect 15160 21916 16344 21944
rect 16868 21944 16896 21975
rect 17034 21972 17040 22024
rect 17092 21972 17098 22024
rect 17126 21972 17132 22024
rect 17184 22012 17190 22024
rect 17497 22015 17555 22021
rect 17497 22012 17509 22015
rect 17184 21984 17509 22012
rect 17184 21972 17190 21984
rect 17497 21981 17509 21984
rect 17543 21981 17555 22015
rect 17497 21975 17555 21981
rect 19242 21972 19248 22024
rect 19300 22012 19306 22024
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 19300 21984 19441 22012
rect 19300 21972 19306 21984
rect 19429 21981 19441 21984
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 19705 22015 19763 22021
rect 19705 21981 19717 22015
rect 19751 21981 19763 22015
rect 19705 21975 19763 21981
rect 16942 21944 16948 21956
rect 16868 21916 16948 21944
rect 15160 21904 15166 21916
rect 16942 21904 16948 21916
rect 17000 21944 17006 21956
rect 19334 21944 19340 21956
rect 17000 21916 19340 21944
rect 17000 21904 17006 21916
rect 17604 21888 17632 21916
rect 19334 21904 19340 21916
rect 19392 21904 19398 21956
rect 19720 21944 19748 21975
rect 19444 21916 19748 21944
rect 19444 21888 19472 21916
rect 3989 21879 4047 21885
rect 3989 21876 4001 21879
rect 3896 21848 4001 21876
rect 3989 21845 4001 21848
rect 4035 21845 4047 21879
rect 3989 21839 4047 21845
rect 4338 21836 4344 21888
rect 4396 21836 4402 21888
rect 5810 21836 5816 21888
rect 5868 21836 5874 21888
rect 6914 21836 6920 21888
rect 6972 21876 6978 21888
rect 8110 21876 8116 21888
rect 6972 21848 8116 21876
rect 6972 21836 6978 21848
rect 8110 21836 8116 21848
rect 8168 21876 8174 21888
rect 8205 21879 8263 21885
rect 8205 21876 8217 21879
rect 8168 21848 8217 21876
rect 8168 21836 8174 21848
rect 8205 21845 8217 21848
rect 8251 21845 8263 21879
rect 8205 21839 8263 21845
rect 8478 21836 8484 21888
rect 8536 21876 8542 21888
rect 9401 21879 9459 21885
rect 9401 21876 9413 21879
rect 8536 21848 9413 21876
rect 8536 21836 8542 21848
rect 9401 21845 9413 21848
rect 9447 21845 9459 21879
rect 9401 21839 9459 21845
rect 9766 21836 9772 21888
rect 9824 21836 9830 21888
rect 9861 21879 9919 21885
rect 9861 21845 9873 21879
rect 9907 21876 9919 21879
rect 10870 21876 10876 21888
rect 9907 21848 10876 21876
rect 9907 21845 9919 21848
rect 9861 21839 9919 21845
rect 10870 21836 10876 21848
rect 10928 21836 10934 21888
rect 11698 21836 11704 21888
rect 11756 21836 11762 21888
rect 11790 21836 11796 21888
rect 11848 21836 11854 21888
rect 12158 21836 12164 21888
rect 12216 21876 12222 21888
rect 12529 21879 12587 21885
rect 12529 21876 12541 21879
rect 12216 21848 12541 21876
rect 12216 21836 12222 21848
rect 12529 21845 12541 21848
rect 12575 21845 12587 21879
rect 12529 21839 12587 21845
rect 12621 21879 12679 21885
rect 12621 21845 12633 21879
rect 12667 21876 12679 21879
rect 12986 21876 12992 21888
rect 12667 21848 12992 21876
rect 12667 21845 12679 21848
rect 12621 21839 12679 21845
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 16206 21836 16212 21888
rect 16264 21876 16270 21888
rect 16761 21879 16819 21885
rect 16761 21876 16773 21879
rect 16264 21848 16773 21876
rect 16264 21836 16270 21848
rect 16761 21845 16773 21848
rect 16807 21845 16819 21879
rect 16761 21839 16819 21845
rect 17586 21836 17592 21888
rect 17644 21836 17650 21888
rect 19426 21836 19432 21888
rect 19484 21836 19490 21888
rect 19812 21876 19840 22052
rect 22204 22052 23612 22080
rect 19978 21972 19984 22024
rect 20036 21972 20042 22024
rect 20162 21972 20168 22024
rect 20220 21972 20226 22024
rect 22002 21972 22008 22024
rect 22060 22012 22066 22024
rect 22204 22021 22232 22052
rect 22189 22015 22247 22021
rect 22189 22012 22201 22015
rect 22060 21984 22201 22012
rect 22060 21972 22066 21984
rect 22189 21981 22201 21984
rect 22235 21981 22247 22015
rect 22189 21975 22247 21981
rect 22278 21972 22284 22024
rect 22336 22012 22342 22024
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 22336 21984 22385 22012
rect 22336 21972 22342 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 22741 22015 22799 22021
rect 22741 21981 22753 22015
rect 22787 22012 22799 22015
rect 22925 22015 22983 22021
rect 22925 22012 22937 22015
rect 22787 21984 22937 22012
rect 22787 21981 22799 21984
rect 22741 21975 22799 21981
rect 22925 21981 22937 21984
rect 22971 22012 22983 22015
rect 23474 22012 23480 22024
rect 22971 21984 23480 22012
rect 22971 21981 22983 21984
rect 22925 21975 22983 21981
rect 23474 21972 23480 21984
rect 23532 21972 23538 22024
rect 23584 22021 23612 22052
rect 23661 22049 23673 22083
rect 23707 22080 23719 22083
rect 24026 22080 24032 22092
rect 23707 22052 24032 22080
rect 23707 22049 23719 22052
rect 23661 22043 23719 22049
rect 24026 22040 24032 22052
rect 24084 22040 24090 22092
rect 24964 22080 24992 22108
rect 24964 22052 25084 22080
rect 23569 22015 23627 22021
rect 23569 21981 23581 22015
rect 23615 21981 23627 22015
rect 23569 21975 23627 21981
rect 24486 21972 24492 22024
rect 24544 22012 24550 22024
rect 24673 22015 24731 22021
rect 24673 22012 24685 22015
rect 24544 21984 24685 22012
rect 24544 21972 24550 21984
rect 24673 21981 24685 21984
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 24762 21972 24768 22024
rect 24820 22012 24826 22024
rect 25056 22021 25084 22052
rect 25314 22040 25320 22092
rect 25372 22040 25378 22092
rect 26050 22040 26056 22092
rect 26108 22080 26114 22092
rect 26108 22052 26280 22080
rect 26108 22040 26114 22052
rect 26252 22024 26280 22052
rect 26602 22040 26608 22092
rect 26660 22080 26666 22092
rect 27249 22083 27307 22089
rect 27249 22080 27261 22083
rect 26660 22052 27261 22080
rect 26660 22040 26666 22052
rect 27249 22049 27261 22052
rect 27295 22049 27307 22083
rect 27249 22043 27307 22049
rect 24857 22015 24915 22021
rect 24857 22012 24869 22015
rect 24820 21984 24869 22012
rect 24820 21972 24826 21984
rect 24857 21981 24869 21984
rect 24903 21981 24915 22015
rect 24857 21975 24915 21981
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 21981 25007 22015
rect 24949 21975 25007 21981
rect 25041 22015 25099 22021
rect 25041 21981 25053 22015
rect 25087 21981 25099 22015
rect 25041 21975 25099 21981
rect 19886 21904 19892 21956
rect 19944 21944 19950 21956
rect 20346 21944 20352 21956
rect 19944 21916 20352 21944
rect 19944 21904 19950 21916
rect 20346 21904 20352 21916
rect 20404 21904 20410 21956
rect 22649 21947 22707 21953
rect 22649 21913 22661 21947
rect 22695 21944 22707 21947
rect 23014 21944 23020 21956
rect 22695 21916 23020 21944
rect 22695 21913 22707 21916
rect 22649 21907 22707 21913
rect 23014 21904 23020 21916
rect 23072 21904 23078 21956
rect 23382 21904 23388 21956
rect 23440 21944 23446 21956
rect 24964 21944 24992 21975
rect 25682 21972 25688 22024
rect 25740 21972 25746 22024
rect 25774 21972 25780 22024
rect 25832 21972 25838 22024
rect 26234 22021 26240 22024
rect 26197 22015 26240 22021
rect 26197 21981 26209 22015
rect 26197 21975 26240 21981
rect 26234 21972 26240 21975
rect 26292 21972 26298 22024
rect 26510 21972 26516 22024
rect 26568 22012 26574 22024
rect 27448 22021 27476 22120
rect 27801 22117 27813 22120
rect 27847 22117 27859 22151
rect 28184 22148 28212 22188
rect 28258 22176 28264 22228
rect 28316 22216 28322 22228
rect 28442 22216 28448 22228
rect 28316 22188 28448 22216
rect 28316 22176 28322 22188
rect 28442 22176 28448 22188
rect 28500 22216 28506 22228
rect 32861 22219 32919 22225
rect 32861 22216 32873 22219
rect 28500 22188 28948 22216
rect 28500 22176 28506 22188
rect 28184 22120 28856 22148
rect 27801 22111 27859 22117
rect 27522 22040 27528 22092
rect 27580 22080 27586 22092
rect 27580 22052 28672 22080
rect 27580 22040 27586 22052
rect 28000 22021 28028 22052
rect 27433 22015 27491 22021
rect 27433 22012 27445 22015
rect 26568 21984 27445 22012
rect 26568 21972 26574 21984
rect 27433 21981 27445 21984
rect 27479 21981 27491 22015
rect 27433 21975 27491 21981
rect 27709 22015 27767 22021
rect 27709 21981 27721 22015
rect 27755 21981 27767 22015
rect 27709 21975 27767 21981
rect 27985 22015 28043 22021
rect 27985 21981 27997 22015
rect 28031 21981 28043 22015
rect 27985 21975 28043 21981
rect 28353 22015 28411 22021
rect 28353 21981 28365 22015
rect 28399 22012 28411 22015
rect 28442 22012 28448 22024
rect 28399 21984 28448 22012
rect 28399 21981 28411 21984
rect 28353 21975 28411 21981
rect 23440 21916 24992 21944
rect 25700 21944 25728 21972
rect 25961 21947 26019 21953
rect 25961 21944 25973 21947
rect 25700 21916 25973 21944
rect 23440 21904 23446 21916
rect 25961 21913 25973 21916
rect 26007 21913 26019 21947
rect 25961 21907 26019 21913
rect 26053 21947 26111 21953
rect 26053 21913 26065 21947
rect 26099 21913 26111 21947
rect 26053 21907 26111 21913
rect 22094 21876 22100 21888
rect 19812 21848 22100 21876
rect 22094 21836 22100 21848
rect 22152 21836 22158 21888
rect 22462 21836 22468 21888
rect 22520 21876 22526 21888
rect 26068 21876 26096 21907
rect 27724 21888 27752 21975
rect 28442 21972 28448 21984
rect 28500 21972 28506 22024
rect 28644 22021 28672 22052
rect 28629 22015 28687 22021
rect 28629 21981 28641 22015
rect 28675 21981 28687 22015
rect 28629 21975 28687 21981
rect 28718 21972 28724 22024
rect 28776 22012 28782 22024
rect 28828 22021 28856 22120
rect 28920 22021 28948 22188
rect 31404 22188 32873 22216
rect 30745 22151 30803 22157
rect 30745 22148 30757 22151
rect 30485 22120 30757 22148
rect 30006 22040 30012 22092
rect 30064 22080 30070 22092
rect 30377 22083 30435 22089
rect 30377 22080 30389 22083
rect 30064 22052 30389 22080
rect 30064 22040 30070 22052
rect 30377 22049 30389 22052
rect 30423 22049 30435 22083
rect 30377 22043 30435 22049
rect 28813 22015 28871 22021
rect 28813 22012 28825 22015
rect 28776 21984 28825 22012
rect 28776 21972 28782 21984
rect 28813 21981 28825 21984
rect 28859 21981 28871 22015
rect 28813 21975 28871 21981
rect 28905 22015 28963 22021
rect 28905 21981 28917 22015
rect 28951 21981 28963 22015
rect 28905 21975 28963 21981
rect 28997 22015 29055 22021
rect 28997 21981 29009 22015
rect 29043 22012 29055 22015
rect 29086 22012 29092 22024
rect 29043 21984 29092 22012
rect 29043 21981 29055 21984
rect 28997 21975 29055 21981
rect 29086 21972 29092 21984
rect 29144 21972 29150 22024
rect 30485 21984 30513 22120
rect 30745 22117 30757 22120
rect 30791 22117 30803 22151
rect 30745 22111 30803 22117
rect 31018 22108 31024 22160
rect 31076 22148 31082 22160
rect 31076 22120 31340 22148
rect 31076 22108 31082 22120
rect 31312 22089 31340 22120
rect 31297 22083 31355 22089
rect 31297 22049 31309 22083
rect 31343 22049 31355 22083
rect 31297 22043 31355 22049
rect 30558 21972 30564 22024
rect 30616 22012 30622 22024
rect 31205 22015 31263 22021
rect 31205 22012 31217 22015
rect 30616 21984 31217 22012
rect 30616 21972 30622 21984
rect 31205 21981 31217 21984
rect 31251 22012 31263 22015
rect 31404 22012 31432 22188
rect 32861 22185 32873 22188
rect 32907 22185 32919 22219
rect 33226 22216 33232 22228
rect 32861 22179 32919 22185
rect 33066 22188 33232 22216
rect 31938 22108 31944 22160
rect 31996 22148 32002 22160
rect 32125 22151 32183 22157
rect 32125 22148 32137 22151
rect 31996 22120 32137 22148
rect 31996 22108 32002 22120
rect 32125 22117 32137 22120
rect 32171 22117 32183 22151
rect 32493 22151 32551 22157
rect 32493 22148 32505 22151
rect 32125 22111 32183 22117
rect 32232 22120 32505 22148
rect 31251 21984 31432 22012
rect 31251 21981 31263 21984
rect 31205 21975 31263 21981
rect 31846 21972 31852 22024
rect 31904 21972 31910 22024
rect 31941 22015 31999 22021
rect 31941 21981 31953 22015
rect 31987 22012 31999 22015
rect 32030 22012 32036 22024
rect 31987 21984 32036 22012
rect 31987 21981 31999 21984
rect 31941 21975 31999 21981
rect 32030 21972 32036 21984
rect 32088 21972 32094 22024
rect 32125 22015 32183 22021
rect 32125 21981 32137 22015
rect 32171 22012 32183 22015
rect 32232 22012 32260 22120
rect 32493 22117 32505 22120
rect 32539 22148 32551 22151
rect 32766 22148 32772 22160
rect 32539 22120 32772 22148
rect 32539 22117 32551 22120
rect 32493 22111 32551 22117
rect 32766 22108 32772 22120
rect 32824 22148 32830 22160
rect 33066 22148 33094 22188
rect 33226 22176 33232 22188
rect 33284 22176 33290 22228
rect 33318 22176 33324 22228
rect 33376 22176 33382 22228
rect 36170 22216 36176 22228
rect 35728 22188 36176 22216
rect 33336 22148 33364 22176
rect 32824 22120 33094 22148
rect 33152 22120 33364 22148
rect 32824 22108 32830 22120
rect 33152 22089 33180 22120
rect 32585 22083 32643 22089
rect 32585 22049 32597 22083
rect 32631 22080 32643 22083
rect 33137 22083 33195 22089
rect 33137 22080 33149 22083
rect 32631 22052 33149 22080
rect 32631 22049 32643 22052
rect 32585 22043 32643 22049
rect 33137 22049 33149 22052
rect 33183 22049 33195 22083
rect 33137 22043 33195 22049
rect 33226 22040 33232 22092
rect 33284 22040 33290 22092
rect 33321 22083 33379 22089
rect 33321 22049 33333 22083
rect 33367 22080 33379 22083
rect 33502 22080 33508 22092
rect 33367 22052 33508 22080
rect 33367 22049 33379 22052
rect 33321 22043 33379 22049
rect 33502 22040 33508 22052
rect 33560 22040 33566 22092
rect 35345 22083 35403 22089
rect 35345 22049 35357 22083
rect 35391 22080 35403 22083
rect 35618 22080 35624 22092
rect 35391 22052 35624 22080
rect 35391 22049 35403 22052
rect 35345 22043 35403 22049
rect 35618 22040 35624 22052
rect 35676 22040 35682 22092
rect 35728 22089 35756 22188
rect 36170 22176 36176 22188
rect 36228 22176 36234 22228
rect 35912 22120 36216 22148
rect 35713 22083 35771 22089
rect 35713 22049 35725 22083
rect 35759 22049 35771 22083
rect 35713 22043 35771 22049
rect 35805 22083 35863 22089
rect 35805 22049 35817 22083
rect 35851 22080 35863 22083
rect 35912 22080 35940 22120
rect 35851 22052 35940 22080
rect 35989 22083 36047 22089
rect 35851 22049 35863 22052
rect 35805 22043 35863 22049
rect 35989 22049 36001 22083
rect 36035 22080 36047 22083
rect 36078 22080 36084 22092
rect 36035 22052 36084 22080
rect 36035 22049 36047 22052
rect 35989 22043 36047 22049
rect 36078 22040 36084 22052
rect 36136 22040 36142 22092
rect 32171 21984 32260 22012
rect 32401 22015 32459 22021
rect 32171 21981 32183 21984
rect 32125 21975 32183 21981
rect 32401 21981 32413 22015
rect 32447 21981 32459 22015
rect 32401 21975 32459 21981
rect 28169 21947 28227 21953
rect 28169 21944 28181 21947
rect 27816 21916 28181 21944
rect 27816 21888 27844 21916
rect 28169 21913 28181 21916
rect 28215 21913 28227 21947
rect 28169 21907 28227 21913
rect 22520 21848 26096 21876
rect 26346 21879 26404 21885
rect 22520 21836 22526 21848
rect 26346 21845 26358 21879
rect 26392 21876 26404 21879
rect 27522 21876 27528 21888
rect 26392 21848 27528 21876
rect 26392 21845 26404 21848
rect 26346 21839 26404 21845
rect 27522 21836 27528 21848
rect 27580 21836 27586 21888
rect 27614 21836 27620 21888
rect 27672 21836 27678 21888
rect 27706 21836 27712 21888
rect 27764 21836 27770 21888
rect 27798 21836 27804 21888
rect 27856 21836 27862 21888
rect 28184 21876 28212 21907
rect 28258 21904 28264 21956
rect 28316 21904 28322 21956
rect 29825 21947 29883 21953
rect 28368 21916 29776 21944
rect 28368 21876 28396 21916
rect 28184 21848 28396 21876
rect 28534 21836 28540 21888
rect 28592 21836 28598 21888
rect 28994 21836 29000 21888
rect 29052 21876 29058 21888
rect 29181 21879 29239 21885
rect 29181 21876 29193 21879
rect 29052 21848 29193 21876
rect 29052 21836 29058 21848
rect 29181 21845 29193 21848
rect 29227 21845 29239 21879
rect 29748 21876 29776 21916
rect 29825 21913 29837 21947
rect 29871 21944 29883 21947
rect 29871 21916 30512 21944
rect 29871 21913 29883 21916
rect 29825 21907 29883 21913
rect 30484 21888 30512 21916
rect 31110 21904 31116 21956
rect 31168 21944 31174 21956
rect 32217 21947 32275 21953
rect 31168 21916 31754 21944
rect 31168 21904 31174 21916
rect 30374 21876 30380 21888
rect 29748 21848 30380 21876
rect 29181 21839 29239 21845
rect 30374 21836 30380 21848
rect 30432 21836 30438 21888
rect 30466 21836 30472 21888
rect 30524 21836 30530 21888
rect 31726 21876 31754 21916
rect 32217 21913 32229 21947
rect 32263 21913 32275 21947
rect 32416 21944 32444 21975
rect 32674 21972 32680 22024
rect 32732 21972 32738 22024
rect 33045 22015 33103 22021
rect 33045 21981 33057 22015
rect 33091 22012 33103 22015
rect 34422 22012 34428 22024
rect 33091 21984 34428 22012
rect 33091 21981 33103 21984
rect 33045 21975 33103 21981
rect 34422 21972 34428 21984
rect 34480 21972 34486 22024
rect 34790 21972 34796 22024
rect 34848 22012 34854 22024
rect 35069 22015 35127 22021
rect 35069 22012 35081 22015
rect 34848 21984 35081 22012
rect 34848 21972 34854 21984
rect 35069 21981 35081 21984
rect 35115 21981 35127 22015
rect 35069 21975 35127 21981
rect 35250 21972 35256 22024
rect 35308 22012 35314 22024
rect 35897 22015 35955 22021
rect 35897 22012 35909 22015
rect 35308 21984 35909 22012
rect 35308 21972 35314 21984
rect 35897 21981 35909 21984
rect 35943 21981 35955 22015
rect 35897 21975 35955 21981
rect 32582 21944 32588 21956
rect 32416 21916 32588 21944
rect 32217 21907 32275 21913
rect 32232 21876 32260 21907
rect 32582 21904 32588 21916
rect 32640 21904 32646 21956
rect 34440 21944 34468 21972
rect 35161 21947 35219 21953
rect 35161 21944 35173 21947
rect 34440 21916 35173 21944
rect 35161 21913 35173 21916
rect 35207 21913 35219 21947
rect 35161 21907 35219 21913
rect 31726 21848 32260 21876
rect 34698 21836 34704 21888
rect 34756 21836 34762 21888
rect 35176 21876 35204 21907
rect 35529 21879 35587 21885
rect 35529 21876 35541 21879
rect 35176 21848 35541 21876
rect 35529 21845 35541 21848
rect 35575 21845 35587 21879
rect 35529 21839 35587 21845
rect 35710 21836 35716 21888
rect 35768 21876 35774 21888
rect 36188 21876 36216 22120
rect 36446 22040 36452 22092
rect 36504 22080 36510 22092
rect 37001 22083 37059 22089
rect 37001 22080 37013 22083
rect 36504 22052 37013 22080
rect 36504 22040 36510 22052
rect 37001 22049 37013 22052
rect 37047 22049 37059 22083
rect 37001 22043 37059 22049
rect 36817 22015 36875 22021
rect 36817 21981 36829 22015
rect 36863 22012 36875 22015
rect 36906 22012 36912 22024
rect 36863 21984 36912 22012
rect 36863 21981 36875 21984
rect 36817 21975 36875 21981
rect 36906 21972 36912 21984
rect 36964 21972 36970 22024
rect 36633 21879 36691 21885
rect 36633 21876 36645 21879
rect 35768 21848 36645 21876
rect 35768 21836 35774 21848
rect 36633 21845 36645 21848
rect 36679 21845 36691 21879
rect 36633 21839 36691 21845
rect 1104 21786 38272 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38272 21786
rect 1104 21712 38272 21734
rect 1762 21632 1768 21684
rect 1820 21632 1826 21684
rect 1946 21632 1952 21684
rect 2004 21672 2010 21684
rect 3237 21675 3295 21681
rect 3237 21672 3249 21675
rect 2004 21644 3249 21672
rect 2004 21632 2010 21644
rect 3237 21641 3249 21644
rect 3283 21641 3295 21675
rect 3237 21635 3295 21641
rect 4338 21632 4344 21684
rect 4396 21632 4402 21684
rect 4706 21672 4712 21684
rect 4540 21644 4712 21672
rect 1673 21607 1731 21613
rect 1673 21573 1685 21607
rect 1719 21604 1731 21607
rect 1780 21604 1808 21632
rect 1719 21576 1808 21604
rect 1719 21573 1731 21576
rect 1673 21567 1731 21573
rect 2774 21496 2780 21548
rect 2832 21496 2838 21548
rect 3602 21536 3608 21548
rect 3160 21508 3608 21536
rect 1394 21428 1400 21480
rect 1452 21428 1458 21480
rect 3160 21477 3188 21508
rect 3602 21496 3608 21508
rect 3660 21496 3666 21548
rect 4356 21545 4384 21632
rect 4540 21613 4568 21644
rect 4706 21632 4712 21644
rect 4764 21632 4770 21684
rect 4908 21644 8340 21672
rect 4540 21607 4609 21613
rect 4540 21576 4563 21607
rect 4551 21573 4563 21576
rect 4597 21573 4609 21607
rect 4551 21567 4609 21573
rect 3697 21539 3755 21545
rect 3697 21505 3709 21539
rect 3743 21536 3755 21539
rect 4065 21539 4123 21545
rect 4065 21536 4077 21539
rect 3743 21508 4077 21536
rect 3743 21505 3755 21508
rect 3697 21499 3755 21505
rect 4065 21505 4077 21508
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 4249 21539 4307 21545
rect 4249 21505 4261 21539
rect 4295 21505 4307 21539
rect 4249 21499 4307 21505
rect 4341 21539 4399 21545
rect 4341 21505 4353 21539
rect 4387 21505 4399 21539
rect 4341 21499 4399 21505
rect 4433 21539 4491 21545
rect 4433 21505 4445 21539
rect 4479 21505 4491 21539
rect 4433 21499 4491 21505
rect 4709 21539 4767 21545
rect 4709 21505 4721 21539
rect 4755 21536 4767 21539
rect 4908 21536 4936 21644
rect 5166 21564 5172 21616
rect 5224 21564 5230 21616
rect 6914 21604 6920 21616
rect 5276 21576 6920 21604
rect 4755 21508 4936 21536
rect 4985 21539 5043 21545
rect 4755 21505 4767 21508
rect 4709 21499 4767 21505
rect 4985 21505 4997 21539
rect 5031 21536 5043 21539
rect 5276 21536 5304 21576
rect 6914 21564 6920 21576
rect 6972 21564 6978 21616
rect 7282 21564 7288 21616
rect 7340 21564 7346 21616
rect 5031 21508 5304 21536
rect 5031 21505 5043 21508
rect 4985 21499 5043 21505
rect 3145 21471 3203 21477
rect 3145 21437 3157 21471
rect 3191 21437 3203 21471
rect 3145 21431 3203 21437
rect 3881 21471 3939 21477
rect 3881 21437 3893 21471
rect 3927 21437 3939 21471
rect 3881 21431 3939 21437
rect 3050 21292 3056 21344
rect 3108 21332 3114 21344
rect 3896 21332 3924 21431
rect 4264 21400 4292 21499
rect 4448 21468 4476 21499
rect 5718 21496 5724 21548
rect 5776 21496 5782 21548
rect 5810 21496 5816 21548
rect 5868 21496 5874 21548
rect 5905 21539 5963 21545
rect 5905 21505 5917 21539
rect 5951 21505 5963 21539
rect 5905 21499 5963 21505
rect 6089 21539 6147 21545
rect 6089 21505 6101 21539
rect 6135 21536 6147 21539
rect 6178 21536 6184 21548
rect 6135 21508 6184 21536
rect 6135 21505 6147 21508
rect 6089 21499 6147 21505
rect 5353 21471 5411 21477
rect 4448 21440 5120 21468
rect 5092 21412 5120 21440
rect 5353 21437 5365 21471
rect 5399 21468 5411 21471
rect 5920 21468 5948 21499
rect 6178 21496 6184 21508
rect 6236 21496 6242 21548
rect 5399 21440 5948 21468
rect 6549 21471 6607 21477
rect 5399 21437 5411 21440
rect 5353 21431 5411 21437
rect 6549 21437 6561 21471
rect 6595 21468 6607 21471
rect 6595 21440 6684 21468
rect 6595 21437 6607 21440
rect 6549 21431 6607 21437
rect 4614 21400 4620 21412
rect 4264 21372 4620 21400
rect 4614 21360 4620 21372
rect 4672 21360 4678 21412
rect 5074 21360 5080 21412
rect 5132 21360 5138 21412
rect 6656 21344 6684 21440
rect 6822 21428 6828 21480
rect 6880 21428 6886 21480
rect 8312 21412 8340 21644
rect 8846 21632 8852 21684
rect 8904 21672 8910 21684
rect 9125 21675 9183 21681
rect 9125 21672 9137 21675
rect 8904 21644 9137 21672
rect 8904 21632 8910 21644
rect 9125 21641 9137 21644
rect 9171 21641 9183 21675
rect 9125 21635 9183 21641
rect 9306 21632 9312 21684
rect 9364 21672 9370 21684
rect 9769 21675 9827 21681
rect 9769 21672 9781 21675
rect 9364 21644 9781 21672
rect 9364 21632 9370 21644
rect 9769 21641 9781 21644
rect 9815 21641 9827 21675
rect 9769 21635 9827 21641
rect 11238 21632 11244 21684
rect 11296 21672 11302 21684
rect 11517 21675 11575 21681
rect 11517 21672 11529 21675
rect 11296 21644 11529 21672
rect 11296 21632 11302 21644
rect 11517 21641 11529 21644
rect 11563 21641 11575 21675
rect 11517 21635 11575 21641
rect 11885 21675 11943 21681
rect 11885 21641 11897 21675
rect 11931 21672 11943 21675
rect 14734 21672 14740 21684
rect 11931 21644 14740 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 14734 21632 14740 21644
rect 14792 21632 14798 21684
rect 14918 21632 14924 21684
rect 14976 21632 14982 21684
rect 17126 21672 17132 21684
rect 15028 21644 17132 21672
rect 13817 21607 13875 21613
rect 9324 21576 13584 21604
rect 8570 21496 8576 21548
rect 8628 21496 8634 21548
rect 9324 21545 9352 21576
rect 9968 21548 9996 21576
rect 9309 21539 9367 21545
rect 9309 21505 9321 21539
rect 9355 21505 9367 21539
rect 9309 21499 9367 21505
rect 9401 21539 9459 21545
rect 9401 21505 9413 21539
rect 9447 21505 9459 21539
rect 9401 21499 9459 21505
rect 9493 21539 9551 21545
rect 9493 21505 9505 21539
rect 9539 21505 9551 21539
rect 9493 21499 9551 21505
rect 8588 21468 8616 21496
rect 9416 21468 9444 21499
rect 8588 21440 9444 21468
rect 9508 21468 9536 21499
rect 9674 21496 9680 21548
rect 9732 21496 9738 21548
rect 9858 21496 9864 21548
rect 9916 21496 9922 21548
rect 9950 21496 9956 21548
rect 10008 21496 10014 21548
rect 10042 21496 10048 21548
rect 10100 21496 10106 21548
rect 10137 21539 10195 21545
rect 10137 21505 10149 21539
rect 10183 21505 10195 21539
rect 10137 21499 10195 21505
rect 9876 21468 9904 21496
rect 10152 21468 10180 21499
rect 10318 21496 10324 21548
rect 10376 21496 10382 21548
rect 12434 21496 12440 21548
rect 12492 21536 12498 21548
rect 12989 21539 13047 21545
rect 12989 21536 13001 21539
rect 12492 21508 13001 21536
rect 12492 21496 12498 21508
rect 12989 21505 13001 21508
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21536 13323 21539
rect 13354 21536 13360 21548
rect 13311 21508 13360 21536
rect 13311 21505 13323 21508
rect 13265 21499 13323 21505
rect 13354 21496 13360 21508
rect 13412 21496 13418 21548
rect 13556 21545 13584 21576
rect 13817 21573 13829 21607
rect 13863 21604 13875 21607
rect 13906 21604 13912 21616
rect 13863 21576 13912 21604
rect 13863 21573 13875 21576
rect 13817 21567 13875 21573
rect 13906 21564 13912 21576
rect 13964 21564 13970 21616
rect 13998 21564 14004 21616
rect 14056 21604 14062 21616
rect 14056 21576 14596 21604
rect 14056 21564 14062 21576
rect 13541 21539 13599 21545
rect 13541 21505 13553 21539
rect 13587 21536 13599 21539
rect 14090 21536 14096 21548
rect 13587 21508 14096 21536
rect 13587 21505 13599 21508
rect 13541 21499 13599 21505
rect 14090 21496 14096 21508
rect 14148 21496 14154 21548
rect 14182 21496 14188 21548
rect 14240 21536 14246 21548
rect 14277 21539 14335 21545
rect 14277 21536 14289 21539
rect 14240 21508 14289 21536
rect 14240 21496 14246 21508
rect 14277 21505 14289 21508
rect 14323 21505 14335 21539
rect 14277 21499 14335 21505
rect 9508 21440 10180 21468
rect 11974 21428 11980 21480
rect 12032 21428 12038 21480
rect 12158 21428 12164 21480
rect 12216 21428 12222 21480
rect 13630 21428 13636 21480
rect 13688 21428 13694 21480
rect 14292 21468 14320 21499
rect 14366 21496 14372 21548
rect 14424 21536 14430 21548
rect 14568 21545 14596 21576
rect 14461 21539 14519 21545
rect 14461 21536 14473 21539
rect 14424 21508 14473 21536
rect 14424 21496 14430 21508
rect 14461 21505 14473 21508
rect 14507 21505 14519 21539
rect 14461 21499 14519 21505
rect 14553 21539 14611 21545
rect 14553 21505 14565 21539
rect 14599 21536 14611 21539
rect 15028 21536 15056 21644
rect 17126 21632 17132 21644
rect 17184 21632 17190 21684
rect 17313 21675 17371 21681
rect 17313 21641 17325 21675
rect 17359 21672 17371 21675
rect 17402 21672 17408 21684
rect 17359 21644 17408 21672
rect 17359 21641 17371 21644
rect 17313 21635 17371 21641
rect 17402 21632 17408 21644
rect 17460 21632 17466 21684
rect 17494 21632 17500 21684
rect 17552 21672 17558 21684
rect 17681 21675 17739 21681
rect 17681 21672 17693 21675
rect 17552 21644 17693 21672
rect 17552 21632 17558 21644
rect 17681 21641 17693 21644
rect 17727 21641 17739 21675
rect 17681 21635 17739 21641
rect 18966 21632 18972 21684
rect 19024 21632 19030 21684
rect 20070 21672 20076 21684
rect 19076 21644 20076 21672
rect 15930 21604 15936 21616
rect 15115 21576 15424 21604
rect 15115 21545 15143 21576
rect 15396 21548 15424 21576
rect 15487 21576 15936 21604
rect 14599 21508 15056 21536
rect 15100 21539 15158 21545
rect 14599 21505 14611 21508
rect 14553 21499 14611 21505
rect 15100 21505 15112 21539
rect 15146 21505 15158 21539
rect 15100 21499 15158 21505
rect 15194 21496 15200 21548
rect 15252 21496 15258 21548
rect 15286 21496 15292 21548
rect 15344 21496 15350 21548
rect 15378 21496 15384 21548
rect 15436 21496 15442 21548
rect 15487 21545 15515 21576
rect 15930 21564 15936 21576
rect 15988 21604 15994 21616
rect 16298 21604 16304 21616
rect 15988 21576 16304 21604
rect 15988 21564 15994 21576
rect 16298 21564 16304 21576
rect 16356 21564 16362 21616
rect 16574 21564 16580 21616
rect 16632 21604 16638 21616
rect 19076 21604 19104 21644
rect 20070 21632 20076 21644
rect 20128 21632 20134 21684
rect 20162 21632 20168 21684
rect 20220 21632 20226 21684
rect 20346 21632 20352 21684
rect 20404 21632 20410 21684
rect 22186 21632 22192 21684
rect 22244 21672 22250 21684
rect 22925 21675 22983 21681
rect 22925 21672 22937 21675
rect 22244 21644 22937 21672
rect 22244 21632 22250 21644
rect 22925 21641 22937 21644
rect 22971 21641 22983 21675
rect 22925 21635 22983 21641
rect 23569 21675 23627 21681
rect 23569 21641 23581 21675
rect 23615 21672 23627 21675
rect 24670 21672 24676 21684
rect 23615 21644 24676 21672
rect 23615 21641 23627 21644
rect 23569 21635 23627 21641
rect 24670 21632 24676 21644
rect 24728 21632 24734 21684
rect 25130 21672 25136 21684
rect 24964 21644 25136 21672
rect 16632 21576 19104 21604
rect 16632 21564 16638 21576
rect 19334 21564 19340 21616
rect 19392 21604 19398 21616
rect 20180 21604 20208 21632
rect 20364 21604 20392 21632
rect 21174 21604 21180 21616
rect 19392 21576 19840 21604
rect 19392 21564 19398 21576
rect 15472 21539 15530 21545
rect 15472 21505 15484 21539
rect 15518 21505 15530 21539
rect 15472 21499 15530 21505
rect 15565 21539 15623 21545
rect 15565 21505 15577 21539
rect 15611 21536 15623 21539
rect 16942 21536 16948 21548
rect 15611 21508 16948 21536
rect 15611 21505 15623 21508
rect 15565 21499 15623 21505
rect 16942 21496 16948 21508
rect 17000 21496 17006 21548
rect 17126 21496 17132 21548
rect 17184 21536 17190 21548
rect 17497 21539 17555 21545
rect 17497 21536 17509 21539
rect 17184 21508 17509 21536
rect 17184 21496 17190 21508
rect 17497 21505 17509 21508
rect 17543 21505 17555 21539
rect 17497 21499 17555 21505
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 17865 21539 17923 21545
rect 17865 21536 17877 21539
rect 17819 21508 17877 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 17865 21505 17877 21508
rect 17911 21505 17923 21539
rect 17865 21499 17923 21505
rect 17954 21496 17960 21548
rect 18012 21536 18018 21548
rect 19242 21536 19248 21548
rect 18012 21508 19248 21536
rect 18012 21496 18018 21508
rect 19242 21496 19248 21508
rect 19300 21536 19306 21548
rect 19521 21539 19579 21545
rect 19521 21536 19533 21539
rect 19300 21508 19533 21536
rect 19300 21496 19306 21508
rect 19521 21505 19533 21508
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 18046 21468 18052 21480
rect 14292 21440 18052 21468
rect 18046 21428 18052 21440
rect 18104 21428 18110 21480
rect 18138 21428 18144 21480
rect 18196 21428 18202 21480
rect 18509 21471 18567 21477
rect 18509 21437 18521 21471
rect 18555 21468 18567 21471
rect 18966 21468 18972 21480
rect 18555 21440 18972 21468
rect 18555 21437 18567 21440
rect 18509 21431 18567 21437
rect 18966 21428 18972 21440
rect 19024 21428 19030 21480
rect 19426 21428 19432 21480
rect 19484 21428 19490 21480
rect 19812 21477 19840 21576
rect 19904 21576 20208 21604
rect 20272 21576 21180 21604
rect 19904 21545 19932 21576
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21505 19947 21539
rect 19889 21499 19947 21505
rect 20165 21539 20223 21545
rect 20165 21505 20177 21539
rect 20211 21536 20223 21539
rect 20272 21536 20300 21576
rect 21174 21564 21180 21576
rect 21232 21564 21238 21616
rect 22002 21564 22008 21616
rect 22060 21604 22066 21616
rect 23109 21607 23167 21613
rect 23109 21604 23121 21607
rect 22060 21576 23121 21604
rect 22060 21564 22066 21576
rect 23109 21573 23121 21576
rect 23155 21573 23167 21607
rect 23109 21567 23167 21573
rect 23842 21564 23848 21616
rect 23900 21604 23906 21616
rect 24762 21604 24768 21616
rect 23900 21576 24768 21604
rect 23900 21564 23906 21576
rect 24762 21564 24768 21576
rect 24820 21604 24826 21616
rect 24964 21604 24992 21644
rect 25130 21632 25136 21644
rect 25188 21672 25194 21684
rect 26694 21672 26700 21684
rect 25188 21644 26700 21672
rect 25188 21632 25194 21644
rect 26694 21632 26700 21644
rect 26752 21632 26758 21684
rect 27706 21632 27712 21684
rect 27764 21632 27770 21684
rect 29914 21632 29920 21684
rect 29972 21632 29978 21684
rect 30374 21632 30380 21684
rect 30432 21672 30438 21684
rect 32582 21672 32588 21684
rect 30432 21644 32588 21672
rect 30432 21632 30438 21644
rect 32582 21632 32588 21644
rect 32640 21632 32646 21684
rect 33778 21672 33784 21684
rect 33336 21644 33784 21672
rect 24820 21576 24992 21604
rect 25041 21607 25099 21613
rect 24820 21564 24826 21576
rect 25041 21573 25053 21607
rect 25087 21604 25099 21607
rect 25314 21604 25320 21616
rect 25087 21576 25320 21604
rect 25087 21573 25099 21576
rect 25041 21567 25099 21573
rect 25314 21564 25320 21576
rect 25372 21604 25378 21616
rect 25593 21607 25651 21613
rect 25593 21604 25605 21607
rect 25372 21576 25605 21604
rect 25372 21564 25378 21576
rect 25593 21573 25605 21576
rect 25639 21573 25651 21607
rect 25593 21567 25651 21573
rect 25866 21564 25872 21616
rect 25924 21564 25930 21616
rect 27890 21604 27896 21616
rect 27632 21576 27896 21604
rect 20211 21508 20300 21536
rect 20211 21505 20223 21508
rect 20165 21499 20223 21505
rect 20346 21496 20352 21548
rect 20404 21496 20410 21548
rect 23017 21539 23075 21545
rect 23017 21505 23029 21539
rect 23063 21536 23075 21539
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 23063 21508 23397 21536
rect 23063 21505 23075 21508
rect 23017 21499 23075 21505
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 24857 21539 24915 21545
rect 24857 21505 24869 21539
rect 24903 21505 24915 21539
rect 24857 21499 24915 21505
rect 19797 21471 19855 21477
rect 19797 21437 19809 21471
rect 19843 21468 19855 21471
rect 19978 21468 19984 21480
rect 19843 21440 19984 21468
rect 19843 21437 19855 21440
rect 19797 21431 19855 21437
rect 19978 21428 19984 21440
rect 20036 21428 20042 21480
rect 23201 21471 23259 21477
rect 23201 21437 23213 21471
rect 23247 21437 23259 21471
rect 23201 21431 23259 21437
rect 8294 21360 8300 21412
rect 8352 21400 8358 21412
rect 16574 21400 16580 21412
rect 8352 21372 16580 21400
rect 8352 21360 8358 21372
rect 16574 21360 16580 21372
rect 16632 21360 16638 21412
rect 22922 21400 22928 21412
rect 16868 21372 22928 21400
rect 3108 21304 3924 21332
rect 3108 21292 3114 21304
rect 4890 21292 4896 21344
rect 4948 21332 4954 21344
rect 5445 21335 5503 21341
rect 5445 21332 5457 21335
rect 4948 21304 5457 21332
rect 4948 21292 4954 21304
rect 5445 21301 5457 21304
rect 5491 21301 5503 21335
rect 5445 21295 5503 21301
rect 6638 21292 6644 21344
rect 6696 21292 6702 21344
rect 8110 21292 8116 21344
rect 8168 21332 8174 21344
rect 10962 21332 10968 21344
rect 8168 21304 10968 21332
rect 8168 21292 8174 21304
rect 10962 21292 10968 21304
rect 11020 21332 11026 21344
rect 16868 21332 16896 21372
rect 22922 21360 22928 21372
rect 22980 21360 22986 21412
rect 23216 21400 23244 21431
rect 23290 21428 23296 21480
rect 23348 21468 23354 21480
rect 23400 21468 23428 21499
rect 23348 21440 23428 21468
rect 23348 21428 23354 21440
rect 23474 21400 23480 21412
rect 23032 21372 23480 21400
rect 11020 21304 16896 21332
rect 11020 21292 11026 21304
rect 17126 21292 17132 21344
rect 17184 21332 17190 21344
rect 23032 21332 23060 21372
rect 23474 21360 23480 21372
rect 23532 21360 23538 21412
rect 24872 21400 24900 21499
rect 25130 21496 25136 21548
rect 25188 21496 25194 21548
rect 25225 21539 25283 21545
rect 25225 21505 25237 21539
rect 25271 21536 25283 21539
rect 25498 21536 25504 21548
rect 25271 21508 25504 21536
rect 25271 21505 25283 21508
rect 25225 21499 25283 21505
rect 25498 21496 25504 21508
rect 25556 21496 25562 21548
rect 25685 21539 25743 21545
rect 25685 21505 25697 21539
rect 25731 21536 25743 21539
rect 25884 21536 25912 21564
rect 25731 21508 25912 21536
rect 25731 21505 25743 21508
rect 25685 21499 25743 21505
rect 26050 21496 26056 21548
rect 26108 21536 26114 21548
rect 27632 21545 27660 21576
rect 27890 21564 27896 21576
rect 27948 21604 27954 21616
rect 28810 21604 28816 21616
rect 27948 21576 28816 21604
rect 27948 21564 27954 21576
rect 28810 21564 28816 21576
rect 28868 21564 28874 21616
rect 29730 21564 29736 21616
rect 29788 21564 29794 21616
rect 29932 21604 29960 21632
rect 29932 21576 30788 21604
rect 27433 21539 27491 21545
rect 27433 21536 27445 21539
rect 26108 21508 27445 21536
rect 26108 21496 26114 21508
rect 27433 21505 27445 21508
rect 27479 21505 27491 21539
rect 27433 21499 27491 21505
rect 27617 21539 27675 21545
rect 27617 21505 27629 21539
rect 27663 21505 27675 21539
rect 27617 21499 27675 21505
rect 27448 21468 27476 21499
rect 27706 21496 27712 21548
rect 27764 21496 27770 21548
rect 30009 21539 30067 21545
rect 30009 21505 30021 21539
rect 30055 21536 30067 21539
rect 30558 21536 30564 21548
rect 30055 21508 30564 21536
rect 30055 21505 30067 21508
rect 30009 21499 30067 21505
rect 30558 21496 30564 21508
rect 30616 21496 30622 21548
rect 30760 21545 30788 21576
rect 33336 21548 33364 21644
rect 33778 21632 33784 21644
rect 33836 21632 33842 21684
rect 34698 21632 34704 21684
rect 34756 21632 34762 21684
rect 35250 21632 35256 21684
rect 35308 21632 35314 21684
rect 35897 21675 35955 21681
rect 35897 21641 35909 21675
rect 35943 21672 35955 21675
rect 36449 21675 36507 21681
rect 36449 21672 36461 21675
rect 35943 21644 36461 21672
rect 35943 21641 35955 21644
rect 35897 21635 35955 21641
rect 36449 21641 36461 21644
rect 36495 21641 36507 21675
rect 36449 21635 36507 21641
rect 33873 21607 33931 21613
rect 33873 21604 33885 21607
rect 33520 21576 33885 21604
rect 30745 21539 30803 21545
rect 30745 21505 30757 21539
rect 30791 21505 30803 21539
rect 30745 21499 30803 21505
rect 30929 21539 30987 21545
rect 30929 21505 30941 21539
rect 30975 21536 30987 21539
rect 31110 21536 31116 21548
rect 30975 21508 31116 21536
rect 30975 21505 30987 21508
rect 30929 21499 30987 21505
rect 31110 21496 31116 21508
rect 31168 21496 31174 21548
rect 31938 21496 31944 21548
rect 31996 21536 32002 21548
rect 32493 21539 32551 21545
rect 32493 21536 32505 21539
rect 31996 21508 32505 21536
rect 31996 21496 32002 21508
rect 32493 21505 32505 21508
rect 32539 21505 32551 21539
rect 32493 21499 32551 21505
rect 32674 21496 32680 21548
rect 32732 21496 32738 21548
rect 33318 21496 33324 21548
rect 33376 21496 33382 21548
rect 33520 21545 33548 21576
rect 33873 21573 33885 21576
rect 33919 21573 33931 21607
rect 33873 21567 33931 21573
rect 33413 21539 33471 21545
rect 33413 21505 33425 21539
rect 33459 21505 33471 21539
rect 33413 21499 33471 21505
rect 33505 21539 33563 21545
rect 33505 21505 33517 21539
rect 33551 21505 33563 21539
rect 33505 21499 33563 21505
rect 33428 21468 33456 21499
rect 33594 21496 33600 21548
rect 33652 21536 33658 21548
rect 33689 21539 33747 21545
rect 33689 21536 33701 21539
rect 33652 21508 33701 21536
rect 33652 21496 33658 21508
rect 33689 21505 33701 21508
rect 33735 21505 33747 21539
rect 33689 21499 33747 21505
rect 33778 21496 33784 21548
rect 33836 21496 33842 21548
rect 33965 21539 34023 21545
rect 33965 21505 33977 21539
rect 34011 21536 34023 21539
rect 34716 21536 34744 21632
rect 35342 21564 35348 21616
rect 35400 21564 35406 21616
rect 36357 21607 36415 21613
rect 36357 21604 36369 21607
rect 35728 21576 36369 21604
rect 34011 21508 34744 21536
rect 35161 21539 35219 21545
rect 34011 21505 34023 21508
rect 33965 21499 34023 21505
rect 35161 21505 35173 21539
rect 35207 21536 35219 21539
rect 35360 21536 35388 21564
rect 35728 21548 35756 21576
rect 36357 21573 36369 21576
rect 36403 21573 36415 21607
rect 36357 21567 36415 21573
rect 35207 21508 35388 21536
rect 35207 21505 35219 21508
rect 35161 21499 35219 21505
rect 33980 21468 34008 21499
rect 35710 21496 35716 21548
rect 35768 21496 35774 21548
rect 35802 21496 35808 21548
rect 35860 21496 35866 21548
rect 36170 21496 36176 21548
rect 36228 21536 36234 21548
rect 36265 21539 36323 21545
rect 36265 21536 36277 21539
rect 36228 21508 36277 21536
rect 36228 21496 36234 21508
rect 36265 21505 36277 21508
rect 36311 21505 36323 21539
rect 36265 21499 36323 21505
rect 36446 21496 36452 21548
rect 36504 21536 36510 21548
rect 36725 21539 36783 21545
rect 36725 21536 36737 21539
rect 36504 21508 36737 21536
rect 36504 21496 36510 21508
rect 36725 21505 36737 21508
rect 36771 21505 36783 21539
rect 36725 21499 36783 21505
rect 27448 21440 33094 21468
rect 33428 21440 34008 21468
rect 27430 21400 27436 21412
rect 24872 21372 27436 21400
rect 27430 21360 27436 21372
rect 27488 21360 27494 21412
rect 28718 21360 28724 21412
rect 28776 21400 28782 21412
rect 33066 21400 33094 21440
rect 35618 21428 35624 21480
rect 35676 21468 35682 21480
rect 35989 21471 36047 21477
rect 35989 21468 36001 21471
rect 35676 21440 36001 21468
rect 35676 21428 35682 21440
rect 35989 21437 36001 21440
rect 36035 21437 36047 21471
rect 35989 21431 36047 21437
rect 37182 21428 37188 21480
rect 37240 21428 37246 21480
rect 37200 21400 37228 21428
rect 28776 21372 31064 21400
rect 33066 21372 37228 21400
rect 28776 21360 28782 21372
rect 17184 21304 23060 21332
rect 17184 21292 17190 21304
rect 23106 21292 23112 21344
rect 23164 21292 23170 21344
rect 25409 21335 25467 21341
rect 25409 21301 25421 21335
rect 25455 21332 25467 21335
rect 29178 21332 29184 21344
rect 25455 21304 29184 21332
rect 25455 21301 25467 21304
rect 25409 21295 25467 21301
rect 29178 21292 29184 21304
rect 29236 21292 29242 21344
rect 29638 21292 29644 21344
rect 29696 21332 29702 21344
rect 29733 21335 29791 21341
rect 29733 21332 29745 21335
rect 29696 21304 29745 21332
rect 29696 21292 29702 21304
rect 29733 21301 29745 21304
rect 29779 21301 29791 21335
rect 29733 21295 29791 21301
rect 30926 21292 30932 21344
rect 30984 21292 30990 21344
rect 31036 21332 31064 21372
rect 33045 21335 33103 21341
rect 33045 21332 33057 21335
rect 31036 21304 33057 21332
rect 33045 21301 33057 21304
rect 33091 21332 33103 21335
rect 33226 21332 33232 21344
rect 33091 21304 33232 21332
rect 33091 21301 33103 21304
rect 33045 21295 33103 21301
rect 33226 21292 33232 21304
rect 33284 21292 33290 21344
rect 35434 21292 35440 21344
rect 35492 21292 35498 21344
rect 1104 21242 38272 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38272 21242
rect 1104 21168 38272 21190
rect 4341 21131 4399 21137
rect 4341 21097 4353 21131
rect 4387 21128 4399 21131
rect 4614 21128 4620 21140
rect 4387 21100 4620 21128
rect 4387 21097 4399 21100
rect 4341 21091 4399 21097
rect 4614 21088 4620 21100
rect 4672 21088 4678 21140
rect 6822 21088 6828 21140
rect 6880 21128 6886 21140
rect 6917 21131 6975 21137
rect 6917 21128 6929 21131
rect 6880 21100 6929 21128
rect 6880 21088 6886 21100
rect 6917 21097 6929 21100
rect 6963 21097 6975 21131
rect 8294 21128 8300 21140
rect 6917 21091 6975 21097
rect 7668 21100 8300 21128
rect 7193 21063 7251 21069
rect 3528 21032 4200 21060
rect 3528 20936 3556 21032
rect 4062 20952 4068 21004
rect 4120 20952 4126 21004
rect 4172 21001 4200 21032
rect 7193 21029 7205 21063
rect 7239 21029 7251 21063
rect 7193 21023 7251 21029
rect 4157 20995 4215 21001
rect 4157 20961 4169 20995
rect 4203 20961 4215 20995
rect 4157 20955 4215 20961
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 1854 20924 1860 20936
rect 1811 20896 1860 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 3510 20884 3516 20936
rect 3568 20884 3574 20936
rect 3602 20884 3608 20936
rect 3660 20924 3666 20936
rect 3881 20927 3939 20933
rect 3881 20924 3893 20927
rect 3660 20896 3893 20924
rect 3660 20884 3666 20896
rect 3881 20893 3893 20896
rect 3927 20893 3939 20927
rect 3881 20887 3939 20893
rect 3896 20856 3924 20887
rect 3970 20884 3976 20936
rect 4028 20884 4034 20936
rect 5445 20927 5503 20933
rect 5445 20924 5457 20927
rect 4264 20896 5457 20924
rect 4264 20856 4292 20896
rect 5445 20893 5457 20896
rect 5491 20893 5503 20927
rect 6914 20924 6920 20936
rect 5445 20887 5503 20893
rect 5552 20896 6920 20924
rect 3896 20828 4292 20856
rect 5261 20859 5319 20865
rect 5261 20825 5273 20859
rect 5307 20856 5319 20859
rect 5552 20856 5580 20896
rect 6914 20884 6920 20896
rect 6972 20884 6978 20936
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20924 7159 20927
rect 7208 20924 7236 21023
rect 7668 21001 7696 21100
rect 8294 21088 8300 21100
rect 8352 21088 8358 21140
rect 9493 21131 9551 21137
rect 9493 21097 9505 21131
rect 9539 21128 9551 21131
rect 9766 21128 9772 21140
rect 9539 21100 9772 21128
rect 9539 21097 9551 21100
rect 9493 21091 9551 21097
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 10134 21088 10140 21140
rect 10192 21088 10198 21140
rect 12158 21088 12164 21140
rect 12216 21128 12222 21140
rect 14645 21131 14703 21137
rect 12216 21100 14136 21128
rect 12216 21088 12222 21100
rect 13998 21060 14004 21072
rect 8588 21032 10088 21060
rect 7653 20995 7711 21001
rect 7653 20961 7665 20995
rect 7699 20961 7711 20995
rect 7653 20955 7711 20961
rect 7837 20995 7895 21001
rect 7837 20961 7849 20995
rect 7883 20992 7895 20995
rect 7926 20992 7932 21004
rect 7883 20964 7932 20992
rect 7883 20961 7895 20964
rect 7837 20955 7895 20961
rect 7926 20952 7932 20964
rect 7984 20952 7990 21004
rect 7147 20896 7236 20924
rect 7561 20927 7619 20933
rect 7147 20893 7159 20896
rect 7101 20887 7159 20893
rect 7561 20893 7573 20927
rect 7607 20924 7619 20927
rect 8588 20924 8616 21032
rect 10060 21004 10088 21032
rect 12406 21032 14004 21060
rect 12406 21004 12434 21032
rect 13998 21020 14004 21032
rect 14056 21020 14062 21072
rect 14108 21060 14136 21100
rect 14645 21097 14657 21131
rect 14691 21128 14703 21131
rect 14734 21128 14740 21140
rect 14691 21100 14740 21128
rect 14691 21097 14703 21100
rect 14645 21091 14703 21097
rect 14734 21088 14740 21100
rect 14792 21088 14798 21140
rect 15470 21088 15476 21140
rect 15528 21088 15534 21140
rect 16945 21131 17003 21137
rect 16945 21097 16957 21131
rect 16991 21128 17003 21131
rect 17034 21128 17040 21140
rect 16991 21100 17040 21128
rect 16991 21097 17003 21100
rect 16945 21091 17003 21097
rect 17034 21088 17040 21100
rect 17092 21088 17098 21140
rect 17126 21088 17132 21140
rect 17184 21088 17190 21140
rect 18230 21088 18236 21140
rect 18288 21128 18294 21140
rect 18417 21131 18475 21137
rect 18417 21128 18429 21131
rect 18288 21100 18429 21128
rect 18288 21088 18294 21100
rect 18417 21097 18429 21100
rect 18463 21097 18475 21131
rect 18417 21091 18475 21097
rect 18506 21088 18512 21140
rect 18564 21128 18570 21140
rect 18782 21128 18788 21140
rect 18564 21100 18788 21128
rect 18564 21088 18570 21100
rect 18782 21088 18788 21100
rect 18840 21128 18846 21140
rect 18969 21131 19027 21137
rect 18969 21128 18981 21131
rect 18840 21100 18981 21128
rect 18840 21088 18846 21100
rect 18969 21097 18981 21100
rect 19015 21097 19027 21131
rect 20346 21128 20352 21140
rect 18969 21091 19027 21097
rect 20088 21100 20352 21128
rect 15197 21063 15255 21069
rect 15197 21060 15209 21063
rect 14108 21032 15209 21060
rect 15197 21029 15209 21032
rect 15243 21060 15255 21063
rect 17144 21060 17172 21088
rect 15243 21032 17172 21060
rect 15243 21029 15255 21032
rect 15197 21023 15255 21029
rect 17494 21020 17500 21072
rect 17552 21060 17558 21072
rect 20088 21060 20116 21100
rect 20346 21088 20352 21100
rect 20404 21128 20410 21140
rect 21082 21128 21088 21140
rect 20404 21100 21088 21128
rect 20404 21088 20410 21100
rect 21082 21088 21088 21100
rect 21140 21088 21146 21140
rect 21818 21088 21824 21140
rect 21876 21128 21882 21140
rect 25038 21128 25044 21140
rect 21876 21100 25044 21128
rect 21876 21088 21882 21100
rect 25038 21088 25044 21100
rect 25096 21088 25102 21140
rect 25314 21088 25320 21140
rect 25372 21088 25378 21140
rect 26789 21131 26847 21137
rect 26789 21097 26801 21131
rect 26835 21128 26847 21131
rect 26970 21128 26976 21140
rect 26835 21100 26976 21128
rect 26835 21097 26847 21100
rect 26789 21091 26847 21097
rect 26970 21088 26976 21100
rect 27028 21088 27034 21140
rect 27522 21088 27528 21140
rect 27580 21088 27586 21140
rect 30561 21131 30619 21137
rect 30561 21097 30573 21131
rect 30607 21128 30619 21131
rect 30926 21128 30932 21140
rect 30607 21100 30932 21128
rect 30607 21097 30619 21100
rect 30561 21091 30619 21097
rect 30926 21088 30932 21100
rect 30984 21088 30990 21140
rect 33502 21088 33508 21140
rect 33560 21128 33566 21140
rect 35250 21128 35256 21140
rect 33560 21100 35256 21128
rect 33560 21088 33566 21100
rect 35250 21088 35256 21100
rect 35308 21088 35314 21140
rect 35434 21088 35440 21140
rect 35492 21088 35498 21140
rect 21177 21063 21235 21069
rect 17552 21032 20116 21060
rect 20180 21032 21133 21060
rect 17552 21020 17558 21032
rect 9324 20964 9996 20992
rect 7607 20896 8616 20924
rect 7607 20893 7619 20896
rect 7561 20887 7619 20893
rect 8662 20884 8668 20936
rect 8720 20924 8726 20936
rect 9324 20933 9352 20964
rect 9968 20936 9996 20964
rect 10042 20952 10048 21004
rect 10100 20952 10106 21004
rect 12342 20952 12348 21004
rect 12400 20964 12434 21004
rect 20180 20992 20208 21032
rect 14384 20964 20208 20992
rect 20257 20995 20315 21001
rect 12400 20952 12406 20964
rect 8941 20927 8999 20933
rect 8941 20924 8953 20927
rect 8720 20896 8953 20924
rect 8720 20884 8726 20896
rect 8941 20893 8953 20896
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 9582 20884 9588 20936
rect 9640 20884 9646 20936
rect 9950 20884 9956 20936
rect 10008 20884 10014 20936
rect 13906 20884 13912 20936
rect 13964 20924 13970 20936
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 13964 20896 14105 20924
rect 13964 20884 13970 20896
rect 14093 20893 14105 20896
rect 14139 20924 14151 20927
rect 14182 20924 14188 20936
rect 14139 20896 14188 20924
rect 14139 20893 14151 20896
rect 14093 20887 14151 20893
rect 14182 20884 14188 20896
rect 14240 20884 14246 20936
rect 14384 20933 14412 20964
rect 20257 20961 20269 20995
rect 20303 20992 20315 20995
rect 20898 20992 20904 21004
rect 20303 20964 20904 20992
rect 20303 20961 20315 20964
rect 20257 20955 20315 20961
rect 20898 20952 20904 20964
rect 20956 20992 20962 21004
rect 21105 20992 21133 21032
rect 21177 21029 21189 21063
rect 21223 21060 21235 21063
rect 21910 21060 21916 21072
rect 21223 21032 21916 21060
rect 21223 21029 21235 21032
rect 21177 21023 21235 21029
rect 21910 21020 21916 21032
rect 21968 21060 21974 21072
rect 23106 21060 23112 21072
rect 21968 21032 23112 21060
rect 21968 21020 21974 21032
rect 23106 21020 23112 21032
rect 23164 21020 23170 21072
rect 22094 20992 22100 21004
rect 20956 20964 21041 20992
rect 21105 20964 22100 20992
rect 20956 20952 20962 20964
rect 17126 20933 17132 20936
rect 14369 20927 14427 20933
rect 14369 20893 14381 20927
rect 14415 20893 14427 20927
rect 14369 20887 14427 20893
rect 14466 20927 14524 20933
rect 14466 20893 14478 20927
rect 14512 20893 14524 20927
rect 14466 20887 14524 20893
rect 15381 20927 15439 20933
rect 15381 20893 15393 20927
rect 15427 20924 15439 20927
rect 15565 20927 15623 20933
rect 15427 20896 15516 20924
rect 15427 20893 15439 20896
rect 15381 20887 15439 20893
rect 5307 20828 5580 20856
rect 5307 20825 5319 20828
rect 5261 20819 5319 20825
rect 1486 20748 1492 20800
rect 1544 20748 1550 20800
rect 2866 20748 2872 20800
rect 2924 20788 2930 20800
rect 4062 20788 4068 20800
rect 2924 20760 4068 20788
rect 2924 20748 2930 20760
rect 4062 20748 4068 20760
rect 4120 20788 4126 20800
rect 5276 20788 5304 20819
rect 5626 20816 5632 20868
rect 5684 20816 5690 20868
rect 9125 20859 9183 20865
rect 9125 20825 9137 20859
rect 9171 20825 9183 20859
rect 9125 20819 9183 20825
rect 4120 20760 5304 20788
rect 9140 20788 9168 20819
rect 9214 20816 9220 20868
rect 9272 20816 9278 20868
rect 9766 20816 9772 20868
rect 9824 20816 9830 20868
rect 9858 20816 9864 20868
rect 9916 20856 9922 20868
rect 10594 20856 10600 20868
rect 9916 20828 10600 20856
rect 9916 20816 9922 20828
rect 10594 20816 10600 20828
rect 10652 20816 10658 20868
rect 13998 20816 14004 20868
rect 14056 20856 14062 20868
rect 14277 20859 14335 20865
rect 14277 20856 14289 20859
rect 14056 20828 14289 20856
rect 14056 20816 14062 20828
rect 14277 20825 14289 20828
rect 14323 20825 14335 20859
rect 14277 20819 14335 20825
rect 9784 20788 9812 20816
rect 9140 20760 9812 20788
rect 4120 20748 4126 20760
rect 11422 20748 11428 20800
rect 11480 20788 11486 20800
rect 12802 20788 12808 20800
rect 11480 20760 12808 20788
rect 11480 20748 11486 20760
rect 12802 20748 12808 20760
rect 12860 20748 12866 20800
rect 14090 20748 14096 20800
rect 14148 20788 14154 20800
rect 14476 20788 14504 20887
rect 14918 20816 14924 20868
rect 14976 20816 14982 20868
rect 15488 20800 15516 20896
rect 15565 20893 15577 20927
rect 15611 20924 15623 20927
rect 17124 20924 17132 20933
rect 15611 20896 15700 20924
rect 17087 20896 17132 20924
rect 15611 20893 15623 20896
rect 15565 20887 15623 20893
rect 15672 20800 15700 20896
rect 17124 20887 17132 20896
rect 17126 20884 17132 20887
rect 17184 20884 17190 20936
rect 17497 20927 17555 20933
rect 17497 20893 17509 20927
rect 17543 20924 17555 20927
rect 17862 20924 17868 20936
rect 17543 20896 17868 20924
rect 17543 20893 17555 20896
rect 17497 20887 17555 20893
rect 17862 20884 17868 20896
rect 17920 20924 17926 20936
rect 18542 20927 18600 20933
rect 18542 20924 18554 20927
rect 17920 20896 18554 20924
rect 17920 20884 17926 20896
rect 18542 20893 18554 20896
rect 18588 20893 18600 20927
rect 18542 20887 18600 20893
rect 18782 20884 18788 20936
rect 18840 20924 18846 20936
rect 19061 20927 19119 20933
rect 19061 20924 19073 20927
rect 18840 20896 19073 20924
rect 18840 20884 18846 20896
rect 19061 20893 19073 20896
rect 19107 20893 19119 20927
rect 19337 20927 19395 20933
rect 19337 20924 19349 20927
rect 19061 20887 19119 20893
rect 19168 20896 19349 20924
rect 17221 20859 17279 20865
rect 17221 20825 17233 20859
rect 17267 20825 17279 20859
rect 17221 20819 17279 20825
rect 17313 20859 17371 20865
rect 17313 20825 17325 20859
rect 17359 20856 17371 20859
rect 17402 20856 17408 20868
rect 17359 20828 17408 20856
rect 17359 20825 17371 20828
rect 17313 20819 17371 20825
rect 14148 20760 14504 20788
rect 14148 20748 14154 20760
rect 14550 20748 14556 20800
rect 14608 20788 14614 20800
rect 15194 20788 15200 20800
rect 14608 20760 15200 20788
rect 14608 20748 14614 20760
rect 15194 20748 15200 20760
rect 15252 20748 15258 20800
rect 15470 20748 15476 20800
rect 15528 20748 15534 20800
rect 15654 20748 15660 20800
rect 15712 20748 15718 20800
rect 17236 20788 17264 20819
rect 17402 20816 17408 20828
rect 17460 20856 17466 20868
rect 17460 20828 18552 20856
rect 17460 20816 17466 20828
rect 18524 20800 18552 20828
rect 17586 20788 17592 20800
rect 17236 20760 17592 20788
rect 17586 20748 17592 20760
rect 17644 20748 17650 20800
rect 18506 20748 18512 20800
rect 18564 20788 18570 20800
rect 18601 20791 18659 20797
rect 18601 20788 18613 20791
rect 18564 20760 18613 20788
rect 18564 20748 18570 20760
rect 18601 20757 18613 20760
rect 18647 20788 18659 20791
rect 19168 20788 19196 20896
rect 19337 20893 19349 20896
rect 19383 20893 19395 20927
rect 19337 20887 19395 20893
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20924 19579 20927
rect 19978 20924 19984 20936
rect 19567 20896 19984 20924
rect 19567 20893 19579 20896
rect 19521 20887 19579 20893
rect 19978 20884 19984 20896
rect 20036 20884 20042 20936
rect 20165 20927 20223 20933
rect 20165 20893 20177 20927
rect 20211 20893 20223 20927
rect 20165 20887 20223 20893
rect 20180 20856 20208 20887
rect 20346 20884 20352 20936
rect 20404 20884 20410 20936
rect 20438 20884 20444 20936
rect 20496 20924 20502 20936
rect 20533 20927 20591 20933
rect 20533 20924 20545 20927
rect 20496 20896 20545 20924
rect 20496 20884 20502 20896
rect 20533 20893 20545 20896
rect 20579 20893 20591 20927
rect 20533 20887 20591 20893
rect 20626 20927 20684 20933
rect 20626 20893 20638 20927
rect 20672 20893 20684 20927
rect 20626 20887 20684 20893
rect 19352 20828 20208 20856
rect 20364 20856 20392 20884
rect 20641 20856 20669 20887
rect 20806 20884 20812 20936
rect 20864 20884 20870 20936
rect 21013 20933 21041 20964
rect 22094 20952 22100 20964
rect 22152 20952 22158 21004
rect 22922 20992 22928 21004
rect 22480 20964 22928 20992
rect 20998 20927 21056 20933
rect 20998 20893 21010 20927
rect 21044 20893 21056 20927
rect 20998 20887 21056 20893
rect 20364 20828 20669 20856
rect 20901 20859 20959 20865
rect 19352 20800 19380 20828
rect 20901 20825 20913 20859
rect 20947 20825 20959 20859
rect 21013 20856 21041 20887
rect 21174 20884 21180 20936
rect 21232 20924 21238 20936
rect 21361 20927 21419 20933
rect 21361 20924 21373 20927
rect 21232 20896 21373 20924
rect 21232 20884 21238 20896
rect 21361 20893 21373 20896
rect 21407 20893 21419 20927
rect 21361 20887 21419 20893
rect 21450 20884 21456 20936
rect 21508 20884 21514 20936
rect 21818 20884 21824 20936
rect 21876 20933 21882 20936
rect 21876 20887 21884 20933
rect 21876 20884 21882 20887
rect 22186 20884 22192 20936
rect 22244 20884 22250 20936
rect 22370 20884 22376 20936
rect 22428 20884 22434 20936
rect 22480 20933 22508 20964
rect 22922 20952 22928 20964
rect 22980 20992 22986 21004
rect 23382 20992 23388 21004
rect 22980 20964 23388 20992
rect 22980 20952 22986 20964
rect 23382 20952 23388 20964
rect 23440 20952 23446 21004
rect 24946 20952 24952 21004
rect 25004 20992 25010 21004
rect 25133 20995 25191 21001
rect 25133 20992 25145 20995
rect 25004 20964 25145 20992
rect 25004 20952 25010 20964
rect 25133 20961 25145 20964
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 22465 20927 22523 20933
rect 22465 20893 22477 20927
rect 22511 20893 22523 20927
rect 22465 20887 22523 20893
rect 22557 20927 22615 20933
rect 22557 20893 22569 20927
rect 22603 20924 22615 20927
rect 24394 20924 24400 20936
rect 22603 20896 24400 20924
rect 22603 20893 22615 20896
rect 22557 20887 22615 20893
rect 24394 20884 24400 20896
rect 24452 20884 24458 20936
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 25332 20933 25360 21088
rect 25498 21020 25504 21072
rect 25556 21060 25562 21072
rect 25682 21060 25688 21072
rect 25556 21032 25688 21060
rect 25556 21020 25562 21032
rect 25682 21020 25688 21032
rect 25740 21020 25746 21072
rect 27540 21060 27568 21088
rect 34330 21060 34336 21072
rect 27540 21032 34336 21060
rect 34330 21020 34336 21032
rect 34388 21020 34394 21072
rect 35342 21060 35348 21072
rect 34992 21032 35348 21060
rect 26712 20964 27108 20992
rect 26712 20936 26740 20964
rect 25041 20927 25099 20933
rect 25041 20924 25053 20927
rect 24912 20896 25053 20924
rect 24912 20884 24918 20896
rect 25041 20893 25053 20896
rect 25087 20893 25099 20927
rect 25041 20887 25099 20893
rect 25317 20927 25375 20933
rect 25317 20893 25329 20927
rect 25363 20893 25375 20927
rect 25317 20887 25375 20893
rect 21637 20859 21695 20865
rect 21637 20856 21649 20859
rect 21013 20828 21649 20856
rect 20901 20819 20959 20825
rect 21637 20825 21649 20828
rect 21683 20825 21695 20859
rect 21637 20819 21695 20825
rect 21729 20859 21787 20865
rect 21729 20825 21741 20859
rect 21775 20825 21787 20859
rect 24486 20856 24492 20868
rect 21729 20819 21787 20825
rect 22756 20828 24492 20856
rect 18647 20760 19196 20788
rect 18647 20757 18659 20760
rect 18601 20751 18659 20757
rect 19334 20748 19340 20800
rect 19392 20748 19398 20800
rect 19429 20791 19487 20797
rect 19429 20757 19441 20791
rect 19475 20788 19487 20791
rect 20346 20788 20352 20800
rect 19475 20760 20352 20788
rect 19475 20757 19487 20760
rect 19429 20751 19487 20757
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 20438 20748 20444 20800
rect 20496 20788 20502 20800
rect 20916 20788 20944 20819
rect 20496 20760 20944 20788
rect 20496 20748 20502 20760
rect 21082 20748 21088 20800
rect 21140 20788 21146 20800
rect 21744 20788 21772 20819
rect 21140 20760 21772 20788
rect 21140 20748 21146 20760
rect 22002 20748 22008 20800
rect 22060 20748 22066 20800
rect 22186 20748 22192 20800
rect 22244 20788 22250 20800
rect 22756 20788 22784 20828
rect 24486 20816 24492 20828
rect 24544 20816 24550 20868
rect 22244 20760 22784 20788
rect 22244 20748 22250 20760
rect 22830 20748 22836 20800
rect 22888 20748 22894 20800
rect 24854 20748 24860 20800
rect 24912 20748 24918 20800
rect 25056 20788 25084 20887
rect 26694 20884 26700 20936
rect 26752 20884 26758 20936
rect 27080 20933 27108 20964
rect 27430 20952 27436 21004
rect 27488 20952 27494 21004
rect 27632 20964 30512 20992
rect 26973 20927 27031 20933
rect 26973 20924 26985 20927
rect 26896 20896 26985 20924
rect 26896 20868 26924 20896
rect 26973 20893 26985 20896
rect 27019 20893 27031 20927
rect 26973 20887 27031 20893
rect 27065 20927 27123 20933
rect 27065 20893 27077 20927
rect 27111 20893 27123 20927
rect 27065 20887 27123 20893
rect 27246 20884 27252 20936
rect 27304 20924 27310 20936
rect 27341 20927 27399 20933
rect 27341 20924 27353 20927
rect 27304 20896 27353 20924
rect 27304 20884 27310 20896
rect 27341 20893 27353 20896
rect 27387 20924 27399 20927
rect 27448 20924 27476 20952
rect 27632 20933 27660 20964
rect 30484 20936 30512 20964
rect 30650 20952 30656 21004
rect 30708 20952 30714 21004
rect 32306 20952 32312 21004
rect 32364 20992 32370 21004
rect 33042 20992 33048 21004
rect 32364 20964 33048 20992
rect 32364 20952 32370 20964
rect 33042 20952 33048 20964
rect 33100 20952 33106 21004
rect 34992 20943 35020 21032
rect 35342 21020 35348 21032
rect 35400 21020 35406 21072
rect 35452 20992 35480 21088
rect 35084 20964 35664 20992
rect 34976 20937 35034 20943
rect 27387 20896 27476 20924
rect 27617 20927 27675 20933
rect 27387 20893 27399 20896
rect 27341 20887 27399 20893
rect 27617 20893 27629 20927
rect 27663 20893 27675 20927
rect 27617 20887 27675 20893
rect 27801 20927 27859 20933
rect 27801 20893 27813 20927
rect 27847 20924 27859 20927
rect 29454 20924 29460 20936
rect 27847 20896 29460 20924
rect 27847 20893 27859 20896
rect 27801 20887 27859 20893
rect 29454 20884 29460 20896
rect 29512 20884 29518 20936
rect 30374 20884 30380 20936
rect 30432 20884 30438 20936
rect 30466 20884 30472 20936
rect 30524 20924 30530 20936
rect 33410 20924 33416 20936
rect 30524 20896 33416 20924
rect 30524 20884 30530 20896
rect 33410 20884 33416 20896
rect 33468 20884 33474 20936
rect 34976 20903 34988 20937
rect 35022 20903 35034 20937
rect 35084 20933 35112 20964
rect 34976 20897 35034 20903
rect 35069 20927 35127 20933
rect 35069 20893 35081 20927
rect 35115 20893 35127 20927
rect 35069 20887 35127 20893
rect 35161 20927 35219 20933
rect 35161 20893 35173 20927
rect 35207 20893 35219 20927
rect 35161 20887 35219 20893
rect 26878 20816 26884 20868
rect 26936 20816 26942 20868
rect 27157 20859 27215 20865
rect 27157 20825 27169 20859
rect 27203 20856 27215 20859
rect 27433 20859 27491 20865
rect 27433 20856 27445 20859
rect 27203 20828 27445 20856
rect 27203 20825 27215 20828
rect 27157 20819 27215 20825
rect 27433 20825 27445 20828
rect 27479 20825 27491 20859
rect 27433 20819 27491 20825
rect 27632 20828 31754 20856
rect 27172 20788 27200 20819
rect 27632 20800 27660 20828
rect 25056 20760 27200 20788
rect 27614 20748 27620 20800
rect 27672 20748 27678 20800
rect 30190 20748 30196 20800
rect 30248 20748 30254 20800
rect 31726 20788 31754 20828
rect 33318 20816 33324 20868
rect 33376 20856 33382 20868
rect 34701 20859 34759 20865
rect 34701 20856 34713 20859
rect 33376 20828 34713 20856
rect 33376 20816 33382 20828
rect 34701 20825 34713 20828
rect 34747 20825 34759 20859
rect 35176 20856 35204 20887
rect 35250 20884 35256 20936
rect 35308 20924 35314 20936
rect 35345 20927 35403 20933
rect 35345 20924 35357 20927
rect 35308 20896 35357 20924
rect 35308 20884 35314 20896
rect 35345 20893 35357 20896
rect 35391 20893 35403 20927
rect 35345 20887 35403 20893
rect 35434 20884 35440 20936
rect 35492 20884 35498 20936
rect 35636 20933 35664 20964
rect 35621 20927 35679 20933
rect 35621 20893 35633 20927
rect 35667 20893 35679 20927
rect 35621 20887 35679 20893
rect 37185 20927 37243 20933
rect 37185 20893 37197 20927
rect 37231 20893 37243 20927
rect 37185 20887 37243 20893
rect 35529 20859 35587 20865
rect 35529 20856 35541 20859
rect 35176 20828 35541 20856
rect 34701 20819 34759 20825
rect 35529 20825 35541 20828
rect 35575 20825 35587 20859
rect 35529 20819 35587 20825
rect 37200 20788 37228 20887
rect 37553 20859 37611 20865
rect 37553 20856 37565 20859
rect 37384 20828 37565 20856
rect 37384 20797 37412 20828
rect 37553 20825 37565 20828
rect 37599 20825 37611 20859
rect 37553 20819 37611 20825
rect 31726 20760 37228 20788
rect 37369 20791 37427 20797
rect 37369 20757 37381 20791
rect 37415 20757 37427 20791
rect 37369 20751 37427 20757
rect 37829 20791 37887 20797
rect 37829 20757 37841 20791
rect 37875 20788 37887 20791
rect 37875 20760 38424 20788
rect 37875 20757 37887 20760
rect 37829 20751 37887 20757
rect 38396 20732 38424 20760
rect 1104 20698 38272 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38272 20698
rect 38378 20680 38384 20732
rect 38436 20680 38442 20732
rect 1104 20624 38272 20646
rect 3697 20587 3755 20593
rect 3697 20553 3709 20587
rect 3743 20584 3755 20587
rect 3878 20584 3884 20596
rect 3743 20556 3884 20584
rect 3743 20553 3755 20556
rect 3697 20547 3755 20553
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20448 2835 20451
rect 3142 20448 3148 20460
rect 2823 20420 3148 20448
rect 2823 20417 2835 20420
rect 2777 20411 2835 20417
rect 3142 20408 3148 20420
rect 3200 20448 3206 20460
rect 3513 20451 3571 20457
rect 3200 20420 3372 20448
rect 3200 20408 3206 20420
rect 2866 20340 2872 20392
rect 2924 20340 2930 20392
rect 3050 20340 3056 20392
rect 3108 20340 3114 20392
rect 3344 20389 3372 20420
rect 3513 20417 3525 20451
rect 3559 20448 3571 20451
rect 3602 20448 3608 20460
rect 3559 20420 3608 20448
rect 3559 20417 3571 20420
rect 3513 20411 3571 20417
rect 3602 20408 3608 20420
rect 3660 20408 3666 20460
rect 3804 20457 3832 20556
rect 3878 20544 3884 20556
rect 3936 20544 3942 20596
rect 7561 20587 7619 20593
rect 7561 20553 7573 20587
rect 7607 20584 7619 20587
rect 13170 20584 13176 20596
rect 7607 20556 13176 20584
rect 7607 20553 7619 20556
rect 7561 20547 7619 20553
rect 13170 20544 13176 20556
rect 13228 20544 13234 20596
rect 14274 20544 14280 20596
rect 14332 20544 14338 20596
rect 14829 20587 14887 20593
rect 14829 20553 14841 20587
rect 14875 20584 14887 20587
rect 15562 20584 15568 20596
rect 14875 20556 15568 20584
rect 14875 20553 14887 20556
rect 14829 20547 14887 20553
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 15654 20544 15660 20596
rect 15712 20584 15718 20596
rect 15712 20556 16068 20584
rect 15712 20544 15718 20556
rect 9766 20476 9772 20528
rect 9824 20516 9830 20528
rect 13998 20516 14004 20528
rect 9824 20488 14004 20516
rect 9824 20476 9830 20488
rect 13998 20476 14004 20488
rect 14056 20476 14062 20528
rect 3789 20451 3847 20457
rect 3789 20417 3801 20451
rect 3835 20417 3847 20451
rect 3789 20411 3847 20417
rect 3970 20408 3976 20460
rect 4028 20408 4034 20460
rect 7653 20451 7711 20457
rect 7653 20417 7665 20451
rect 7699 20448 7711 20451
rect 11701 20451 11759 20457
rect 7699 20420 8432 20448
rect 7699 20417 7711 20420
rect 7653 20411 7711 20417
rect 3329 20383 3387 20389
rect 3329 20349 3341 20383
rect 3375 20380 3387 20383
rect 3988 20380 4016 20408
rect 8404 20392 8432 20420
rect 11701 20417 11713 20451
rect 11747 20448 11759 20451
rect 11974 20448 11980 20460
rect 11747 20420 11980 20448
rect 11747 20417 11759 20420
rect 11701 20411 11759 20417
rect 11974 20408 11980 20420
rect 12032 20448 12038 20460
rect 14292 20448 14320 20544
rect 14642 20476 14648 20528
rect 14700 20476 14706 20528
rect 15102 20476 15108 20528
rect 15160 20516 15166 20528
rect 16040 20516 16068 20556
rect 16114 20544 16120 20596
rect 16172 20584 16178 20596
rect 18598 20584 18604 20596
rect 16172 20556 18604 20584
rect 16172 20544 16178 20556
rect 18598 20544 18604 20556
rect 18656 20584 18662 20596
rect 18785 20587 18843 20593
rect 18785 20584 18797 20587
rect 18656 20556 18797 20584
rect 18656 20544 18662 20556
rect 18785 20553 18797 20556
rect 18831 20553 18843 20587
rect 18785 20547 18843 20553
rect 18874 20544 18880 20596
rect 18932 20584 18938 20596
rect 20165 20587 20223 20593
rect 18932 20556 20116 20584
rect 18932 20544 18938 20556
rect 19797 20519 19855 20525
rect 19797 20516 19809 20519
rect 15160 20488 15608 20516
rect 16040 20488 19809 20516
rect 15160 20476 15166 20488
rect 15580 20460 15608 20488
rect 19797 20485 19809 20488
rect 19843 20485 19855 20519
rect 20088 20516 20116 20556
rect 20165 20553 20177 20587
rect 20211 20584 20223 20587
rect 20438 20584 20444 20596
rect 20211 20556 20444 20584
rect 20211 20553 20223 20556
rect 20165 20547 20223 20553
rect 20438 20544 20444 20556
rect 20496 20544 20502 20596
rect 21082 20544 21088 20596
rect 21140 20584 21146 20596
rect 21269 20587 21327 20593
rect 21140 20556 21220 20584
rect 21140 20544 21146 20556
rect 20533 20519 20591 20525
rect 20088 20488 20484 20516
rect 19797 20479 19855 20485
rect 15473 20451 15531 20457
rect 15473 20448 15485 20451
rect 12032 20420 12434 20448
rect 14292 20420 15485 20448
rect 12032 20408 12038 20420
rect 3375 20352 4016 20380
rect 3375 20349 3387 20352
rect 3329 20343 3387 20349
rect 7374 20340 7380 20392
rect 7432 20380 7438 20392
rect 7745 20383 7803 20389
rect 7745 20380 7757 20383
rect 7432 20352 7757 20380
rect 7432 20340 7438 20352
rect 7745 20349 7757 20352
rect 7791 20380 7803 20383
rect 7926 20380 7932 20392
rect 7791 20352 7932 20380
rect 7791 20349 7803 20352
rect 7745 20343 7803 20349
rect 7926 20340 7932 20352
rect 7984 20340 7990 20392
rect 8386 20340 8392 20392
rect 8444 20340 8450 20392
rect 11606 20340 11612 20392
rect 11664 20340 11670 20392
rect 3786 20272 3792 20324
rect 3844 20312 3850 20324
rect 12250 20312 12256 20324
rect 3844 20284 12256 20312
rect 3844 20272 3850 20284
rect 12250 20272 12256 20284
rect 12308 20272 12314 20324
rect 12406 20312 12434 20420
rect 15473 20417 15485 20420
rect 15519 20417 15531 20451
rect 15473 20411 15531 20417
rect 15562 20408 15568 20460
rect 15620 20408 15626 20460
rect 17770 20448 17776 20460
rect 15856 20420 17776 20448
rect 14277 20383 14335 20389
rect 14277 20349 14289 20383
rect 14323 20380 14335 20383
rect 15102 20380 15108 20392
rect 14323 20352 15108 20380
rect 14323 20349 14335 20352
rect 14277 20343 14335 20349
rect 15102 20340 15108 20352
rect 15160 20380 15166 20392
rect 15856 20380 15884 20420
rect 17770 20408 17776 20420
rect 17828 20408 17834 20460
rect 17954 20408 17960 20460
rect 18012 20448 18018 20460
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 18012 20420 18061 20448
rect 18012 20408 18018 20420
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 18138 20408 18144 20460
rect 18196 20448 18202 20460
rect 18414 20448 18420 20460
rect 18196 20420 18420 20448
rect 18196 20408 18202 20420
rect 18414 20408 18420 20420
rect 18472 20408 18478 20460
rect 18506 20408 18512 20460
rect 18564 20408 18570 20460
rect 18598 20408 18604 20460
rect 18656 20408 18662 20460
rect 19242 20448 19248 20460
rect 18708 20420 19248 20448
rect 15160 20352 15884 20380
rect 15933 20383 15991 20389
rect 15160 20340 15166 20352
rect 15933 20349 15945 20383
rect 15979 20380 15991 20383
rect 16114 20380 16120 20392
rect 15979 20352 16120 20380
rect 15979 20349 15991 20352
rect 15933 20343 15991 20349
rect 16114 20340 16120 20352
rect 16172 20340 16178 20392
rect 16942 20340 16948 20392
rect 17000 20380 17006 20392
rect 17589 20383 17647 20389
rect 17589 20380 17601 20383
rect 17000 20352 17601 20380
rect 17000 20340 17006 20352
rect 17589 20349 17601 20352
rect 17635 20349 17647 20383
rect 18708 20380 18736 20420
rect 19242 20408 19248 20420
rect 19300 20408 19306 20460
rect 19981 20451 20039 20457
rect 19981 20417 19993 20451
rect 20027 20448 20039 20451
rect 20070 20448 20076 20460
rect 20027 20420 20076 20448
rect 20027 20417 20039 20420
rect 19981 20411 20039 20417
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20346 20408 20352 20460
rect 20404 20408 20410 20460
rect 17589 20343 17647 20349
rect 18064 20352 18736 20380
rect 18064 20324 18092 20352
rect 19058 20340 19064 20392
rect 19116 20380 19122 20392
rect 19153 20383 19211 20389
rect 19153 20380 19165 20383
rect 19116 20352 19165 20380
rect 19116 20340 19122 20352
rect 19153 20349 19165 20352
rect 19199 20349 19211 20383
rect 20456 20380 20484 20488
rect 20533 20485 20545 20519
rect 20579 20516 20591 20519
rect 20579 20488 21128 20516
rect 20579 20485 20591 20488
rect 20533 20479 20591 20485
rect 20622 20408 20628 20460
rect 20680 20408 20686 20460
rect 20718 20451 20776 20457
rect 20718 20417 20730 20451
rect 20764 20417 20776 20451
rect 20718 20411 20776 20417
rect 20732 20380 20760 20411
rect 20898 20408 20904 20460
rect 20956 20408 20962 20460
rect 21100 20457 21128 20488
rect 20993 20451 21051 20457
rect 20993 20417 21005 20451
rect 21039 20417 21051 20451
rect 20993 20411 21051 20417
rect 21090 20451 21148 20457
rect 21090 20417 21102 20451
rect 21136 20417 21148 20451
rect 21090 20411 21148 20417
rect 20456 20352 20760 20380
rect 21008 20380 21036 20411
rect 21192 20380 21220 20556
rect 21269 20553 21281 20587
rect 21315 20584 21327 20587
rect 23290 20584 23296 20596
rect 21315 20556 23296 20584
rect 21315 20553 21327 20556
rect 21269 20547 21327 20553
rect 23290 20544 23296 20556
rect 23348 20544 23354 20596
rect 23382 20544 23388 20596
rect 23440 20584 23446 20596
rect 25498 20584 25504 20596
rect 23440 20556 25504 20584
rect 23440 20544 23446 20556
rect 25498 20544 25504 20556
rect 25556 20544 25562 20596
rect 27801 20587 27859 20593
rect 27801 20553 27813 20587
rect 27847 20584 27859 20587
rect 27982 20584 27988 20596
rect 27847 20556 27988 20584
rect 27847 20553 27859 20556
rect 27801 20547 27859 20553
rect 27982 20544 27988 20556
rect 28040 20544 28046 20596
rect 35437 20587 35495 20593
rect 35437 20553 35449 20587
rect 35483 20584 35495 20587
rect 35802 20584 35808 20596
rect 35483 20556 35808 20584
rect 35483 20553 35495 20556
rect 35437 20547 35495 20553
rect 35802 20544 35808 20556
rect 35860 20544 35866 20596
rect 27433 20519 27491 20525
rect 27433 20516 27445 20519
rect 24412 20488 27445 20516
rect 24412 20460 24440 20488
rect 27433 20485 27445 20488
rect 27479 20516 27491 20519
rect 32030 20516 32036 20528
rect 27479 20488 32036 20516
rect 27479 20485 27491 20488
rect 27433 20479 27491 20485
rect 32030 20476 32036 20488
rect 32088 20516 32094 20528
rect 33318 20516 33324 20528
rect 32088 20488 33324 20516
rect 32088 20476 32094 20488
rect 33318 20476 33324 20488
rect 33376 20476 33382 20528
rect 24305 20451 24363 20457
rect 24305 20417 24317 20451
rect 24351 20417 24363 20451
rect 24305 20411 24363 20417
rect 21008 20352 21220 20380
rect 19153 20343 19211 20349
rect 22094 20340 22100 20392
rect 22152 20380 22158 20392
rect 23566 20380 23572 20392
rect 22152 20352 23572 20380
rect 22152 20340 22158 20352
rect 23566 20340 23572 20352
rect 23624 20340 23630 20392
rect 12406 20284 17816 20312
rect 17788 20256 17816 20284
rect 18046 20272 18052 20324
rect 18104 20272 18110 20324
rect 22278 20312 22284 20324
rect 18616 20284 22284 20312
rect 18616 20256 18644 20284
rect 22278 20272 22284 20284
rect 22336 20272 22342 20324
rect 24320 20312 24348 20411
rect 24394 20408 24400 20460
rect 24452 20408 24458 20460
rect 24578 20408 24584 20460
rect 24636 20408 24642 20460
rect 24854 20408 24860 20460
rect 24912 20408 24918 20460
rect 25133 20451 25191 20457
rect 25133 20417 25145 20451
rect 25179 20417 25191 20451
rect 25133 20411 25191 20417
rect 24489 20383 24547 20389
rect 24489 20349 24501 20383
rect 24535 20380 24547 20383
rect 24872 20380 24900 20408
rect 24535 20352 24900 20380
rect 24535 20349 24547 20352
rect 24489 20343 24547 20349
rect 24670 20312 24676 20324
rect 24320 20284 24676 20312
rect 24670 20272 24676 20284
rect 24728 20272 24734 20324
rect 25148 20312 25176 20411
rect 25222 20408 25228 20460
rect 25280 20448 25286 20460
rect 25777 20451 25835 20457
rect 25777 20448 25789 20451
rect 25280 20420 25789 20448
rect 25280 20408 25286 20420
rect 25777 20417 25789 20420
rect 25823 20417 25835 20451
rect 25777 20411 25835 20417
rect 25866 20408 25872 20460
rect 25924 20448 25930 20460
rect 25961 20451 26019 20457
rect 25961 20448 25973 20451
rect 25924 20420 25973 20448
rect 25924 20408 25930 20420
rect 25961 20417 25973 20420
rect 26007 20417 26019 20451
rect 25961 20411 26019 20417
rect 26050 20408 26056 20460
rect 26108 20408 26114 20460
rect 26145 20451 26203 20457
rect 26145 20417 26157 20451
rect 26191 20448 26203 20451
rect 26234 20448 26240 20460
rect 26191 20420 26240 20448
rect 26191 20417 26203 20420
rect 26145 20411 26203 20417
rect 26234 20408 26240 20420
rect 26292 20408 26298 20460
rect 26694 20408 26700 20460
rect 26752 20408 26758 20460
rect 27246 20408 27252 20460
rect 27304 20408 27310 20460
rect 27525 20451 27583 20457
rect 27525 20417 27537 20451
rect 27571 20417 27583 20451
rect 27525 20411 27583 20417
rect 25314 20340 25320 20392
rect 25372 20340 25378 20392
rect 25406 20340 25412 20392
rect 25464 20380 25470 20392
rect 25884 20380 25912 20408
rect 25464 20352 25912 20380
rect 25464 20340 25470 20352
rect 26142 20312 26148 20324
rect 25148 20284 26148 20312
rect 26142 20272 26148 20284
rect 26200 20272 26206 20324
rect 2406 20204 2412 20256
rect 2464 20204 2470 20256
rect 3881 20247 3939 20253
rect 3881 20213 3893 20247
rect 3927 20244 3939 20247
rect 3970 20244 3976 20256
rect 3927 20216 3976 20244
rect 3927 20213 3939 20216
rect 3881 20207 3939 20213
rect 3970 20204 3976 20216
rect 4028 20204 4034 20256
rect 7190 20204 7196 20256
rect 7248 20204 7254 20256
rect 11882 20204 11888 20256
rect 11940 20244 11946 20256
rect 11977 20247 12035 20253
rect 11977 20244 11989 20247
rect 11940 20216 11989 20244
rect 11940 20204 11946 20216
rect 11977 20213 11989 20216
rect 12023 20213 12035 20247
rect 11977 20207 12035 20213
rect 14645 20247 14703 20253
rect 14645 20213 14657 20247
rect 14691 20244 14703 20247
rect 16298 20244 16304 20256
rect 14691 20216 16304 20244
rect 14691 20213 14703 20216
rect 14645 20207 14703 20213
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 17770 20204 17776 20256
rect 17828 20204 17834 20256
rect 18598 20204 18604 20256
rect 18656 20204 18662 20256
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 19429 20247 19487 20253
rect 19429 20244 19441 20247
rect 19392 20216 19441 20244
rect 19392 20204 19398 20216
rect 19429 20213 19441 20216
rect 19475 20213 19487 20247
rect 19429 20207 19487 20213
rect 19705 20247 19763 20253
rect 19705 20213 19717 20247
rect 19751 20244 19763 20247
rect 19886 20244 19892 20256
rect 19751 20216 19892 20244
rect 19751 20213 19763 20216
rect 19705 20207 19763 20213
rect 19886 20204 19892 20216
rect 19944 20244 19950 20256
rect 20162 20244 20168 20256
rect 19944 20216 20168 20244
rect 19944 20204 19950 20216
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 20346 20204 20352 20256
rect 20404 20244 20410 20256
rect 21450 20244 21456 20256
rect 20404 20216 21456 20244
rect 20404 20204 20410 20216
rect 21450 20204 21456 20216
rect 21508 20204 21514 20256
rect 21910 20204 21916 20256
rect 21968 20244 21974 20256
rect 24026 20244 24032 20256
rect 21968 20216 24032 20244
rect 21968 20204 21974 20216
rect 24026 20204 24032 20216
rect 24084 20204 24090 20256
rect 24118 20204 24124 20256
rect 24176 20204 24182 20256
rect 24946 20204 24952 20256
rect 25004 20204 25010 20256
rect 25498 20204 25504 20256
rect 25556 20244 25562 20256
rect 26252 20244 26280 20408
rect 26712 20380 26740 20408
rect 27540 20380 27568 20411
rect 27614 20408 27620 20460
rect 27672 20408 27678 20460
rect 28905 20451 28963 20457
rect 28905 20448 28917 20451
rect 28736 20420 28917 20448
rect 28736 20392 28764 20420
rect 28905 20417 28917 20420
rect 28951 20417 28963 20451
rect 28905 20411 28963 20417
rect 29089 20451 29147 20457
rect 29089 20417 29101 20451
rect 29135 20448 29147 20451
rect 29546 20448 29552 20460
rect 29135 20420 29552 20448
rect 29135 20417 29147 20420
rect 29089 20411 29147 20417
rect 26712 20352 27568 20380
rect 27540 20324 27568 20352
rect 28718 20340 28724 20392
rect 28776 20340 28782 20392
rect 28810 20340 28816 20392
rect 28868 20380 28874 20392
rect 29104 20380 29132 20411
rect 29546 20408 29552 20420
rect 29604 20408 29610 20460
rect 29733 20451 29791 20457
rect 29733 20417 29745 20451
rect 29779 20448 29791 20451
rect 30285 20451 30343 20457
rect 30285 20448 30297 20451
rect 29779 20420 30297 20448
rect 29779 20417 29791 20420
rect 29733 20411 29791 20417
rect 30285 20417 30297 20420
rect 30331 20448 30343 20451
rect 30374 20448 30380 20460
rect 30331 20420 30380 20448
rect 30331 20417 30343 20420
rect 30285 20411 30343 20417
rect 30374 20408 30380 20420
rect 30432 20408 30438 20460
rect 30561 20451 30619 20457
rect 30561 20417 30573 20451
rect 30607 20448 30619 20451
rect 30650 20448 30656 20460
rect 30607 20420 30656 20448
rect 30607 20417 30619 20420
rect 30561 20411 30619 20417
rect 30650 20408 30656 20420
rect 30708 20408 30714 20460
rect 30745 20451 30803 20457
rect 30745 20417 30757 20451
rect 30791 20448 30803 20451
rect 30926 20448 30932 20460
rect 30791 20420 30932 20448
rect 30791 20417 30803 20420
rect 30745 20411 30803 20417
rect 30926 20408 30932 20420
rect 30984 20408 30990 20460
rect 31021 20451 31079 20457
rect 31021 20417 31033 20451
rect 31067 20448 31079 20451
rect 31110 20448 31116 20460
rect 31067 20420 31116 20448
rect 31067 20417 31079 20420
rect 31021 20411 31079 20417
rect 31110 20408 31116 20420
rect 31168 20408 31174 20460
rect 32582 20408 32588 20460
rect 32640 20448 32646 20460
rect 33137 20451 33195 20457
rect 33137 20448 33149 20451
rect 32640 20420 33149 20448
rect 32640 20408 32646 20420
rect 33137 20417 33149 20420
rect 33183 20417 33195 20451
rect 33137 20411 33195 20417
rect 35894 20408 35900 20460
rect 35952 20408 35958 20460
rect 28868 20352 29132 20380
rect 28868 20340 28874 20352
rect 29638 20340 29644 20392
rect 29696 20340 29702 20392
rect 29748 20352 31754 20380
rect 26329 20315 26387 20321
rect 26329 20281 26341 20315
rect 26375 20312 26387 20315
rect 27246 20312 27252 20324
rect 26375 20284 27252 20312
rect 26375 20281 26387 20284
rect 26329 20275 26387 20281
rect 27246 20272 27252 20284
rect 27304 20272 27310 20324
rect 27522 20272 27528 20324
rect 27580 20272 27586 20324
rect 28626 20272 28632 20324
rect 28684 20312 28690 20324
rect 29748 20312 29776 20352
rect 28684 20284 29776 20312
rect 28684 20272 28690 20284
rect 30650 20272 30656 20324
rect 30708 20272 30714 20324
rect 31726 20312 31754 20352
rect 33226 20340 33232 20392
rect 33284 20340 33290 20392
rect 34422 20340 34428 20392
rect 34480 20380 34486 20392
rect 35621 20383 35679 20389
rect 35621 20380 35633 20383
rect 34480 20352 35633 20380
rect 34480 20340 34486 20352
rect 35621 20349 35633 20352
rect 35667 20349 35679 20383
rect 35621 20343 35679 20349
rect 35713 20383 35771 20389
rect 35713 20349 35725 20383
rect 35759 20349 35771 20383
rect 35713 20343 35771 20349
rect 33134 20312 33140 20324
rect 31726 20284 33140 20312
rect 33134 20272 33140 20284
rect 33192 20272 33198 20324
rect 33505 20315 33563 20321
rect 33505 20281 33517 20315
rect 33551 20312 33563 20315
rect 34514 20312 34520 20324
rect 33551 20284 34520 20312
rect 33551 20281 33563 20284
rect 33505 20275 33563 20281
rect 34514 20272 34520 20284
rect 34572 20272 34578 20324
rect 35728 20312 35756 20343
rect 35802 20340 35808 20392
rect 35860 20340 35866 20392
rect 34808 20284 35756 20312
rect 34808 20256 34836 20284
rect 25556 20216 26280 20244
rect 25556 20204 25562 20216
rect 28902 20204 28908 20256
rect 28960 20204 28966 20256
rect 30009 20247 30067 20253
rect 30009 20213 30021 20247
rect 30055 20244 30067 20247
rect 31202 20244 31208 20256
rect 30055 20216 31208 20244
rect 30055 20213 30067 20216
rect 30009 20207 30067 20213
rect 31202 20204 31208 20216
rect 31260 20204 31266 20256
rect 34790 20204 34796 20256
rect 34848 20204 34854 20256
rect 1104 20154 38272 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38272 20154
rect 1104 20080 38272 20102
rect 2406 20000 2412 20052
rect 2464 20000 2470 20052
rect 2866 20000 2872 20052
rect 2924 20040 2930 20052
rect 3789 20043 3847 20049
rect 3789 20040 3801 20043
rect 2924 20012 3801 20040
rect 2924 20000 2930 20012
rect 3789 20009 3801 20012
rect 3835 20009 3847 20043
rect 7466 20040 7472 20052
rect 3789 20003 3847 20009
rect 4448 20012 7472 20040
rect 1949 19839 2007 19845
rect 1949 19805 1961 19839
rect 1995 19836 2007 19839
rect 2424 19836 2452 20000
rect 2961 19907 3019 19913
rect 2961 19873 2973 19907
rect 3007 19873 3019 19907
rect 2961 19867 3019 19873
rect 1995 19808 2452 19836
rect 1995 19805 2007 19808
rect 1949 19799 2007 19805
rect 2976 19712 3004 19867
rect 3050 19864 3056 19916
rect 3108 19904 3114 19916
rect 4448 19913 4476 20012
rect 7466 20000 7472 20012
rect 7524 20040 7530 20052
rect 7524 20012 7972 20040
rect 7524 20000 7530 20012
rect 7944 19984 7972 20012
rect 8110 20000 8116 20052
rect 8168 20040 8174 20052
rect 9769 20043 9827 20049
rect 8168 20012 8524 20040
rect 8168 20000 8174 20012
rect 5077 19975 5135 19981
rect 4540 19944 4936 19972
rect 4433 19907 4491 19913
rect 3108 19876 4384 19904
rect 3108 19864 3114 19876
rect 3329 19839 3387 19845
rect 3329 19805 3341 19839
rect 3375 19836 3387 19839
rect 3786 19836 3792 19848
rect 3375 19808 3792 19836
rect 3375 19805 3387 19808
rect 3329 19799 3387 19805
rect 3786 19796 3792 19808
rect 3844 19796 3850 19848
rect 3878 19796 3884 19848
rect 3936 19836 3942 19848
rect 3973 19839 4031 19845
rect 3973 19836 3985 19839
rect 3936 19808 3985 19836
rect 3936 19796 3942 19808
rect 3973 19805 3985 19808
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19805 4123 19839
rect 4356 19836 4384 19876
rect 4433 19873 4445 19907
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 4540 19836 4568 19944
rect 4798 19864 4804 19916
rect 4856 19864 4862 19916
rect 4908 19904 4936 19944
rect 5077 19941 5089 19975
rect 5123 19972 5135 19975
rect 5123 19944 6408 19972
rect 5123 19941 5135 19944
rect 5077 19935 5135 19941
rect 5721 19907 5779 19913
rect 5721 19904 5733 19907
rect 4908 19876 5733 19904
rect 5721 19873 5733 19876
rect 5767 19873 5779 19907
rect 5721 19867 5779 19873
rect 4356 19808 4568 19836
rect 4709 19839 4767 19845
rect 4065 19799 4123 19805
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 5537 19839 5595 19845
rect 5537 19836 5549 19839
rect 4755 19808 5549 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 5537 19805 5549 19808
rect 5583 19836 5595 19839
rect 5902 19836 5908 19848
rect 5583 19808 5908 19836
rect 5583 19805 5595 19808
rect 5537 19799 5595 19805
rect 4080 19768 4108 19799
rect 5902 19796 5908 19808
rect 5960 19796 5966 19848
rect 6380 19845 6408 19944
rect 7926 19932 7932 19984
rect 7984 19932 7990 19984
rect 8389 19975 8447 19981
rect 8389 19941 8401 19975
rect 8435 19941 8447 19975
rect 8496 19972 8524 20012
rect 9769 20009 9781 20043
rect 9815 20040 9827 20043
rect 10226 20040 10232 20052
rect 9815 20012 10232 20040
rect 9815 20009 9827 20012
rect 9769 20003 9827 20009
rect 10226 20000 10232 20012
rect 10284 20000 10290 20052
rect 11606 20000 11612 20052
rect 11664 20000 11670 20052
rect 13817 20043 13875 20049
rect 13817 20009 13829 20043
rect 13863 20040 13875 20043
rect 13998 20040 14004 20052
rect 13863 20012 14004 20040
rect 13863 20009 13875 20012
rect 13817 20003 13875 20009
rect 13998 20000 14004 20012
rect 14056 20000 14062 20052
rect 14090 20000 14096 20052
rect 14148 20040 14154 20052
rect 14737 20043 14795 20049
rect 14737 20040 14749 20043
rect 14148 20012 14749 20040
rect 14148 20000 14154 20012
rect 14737 20009 14749 20012
rect 14783 20009 14795 20043
rect 14737 20003 14795 20009
rect 15565 20043 15623 20049
rect 15565 20009 15577 20043
rect 15611 20040 15623 20043
rect 16114 20040 16120 20052
rect 15611 20012 16120 20040
rect 15611 20009 15623 20012
rect 15565 20003 15623 20009
rect 10413 19975 10471 19981
rect 8496 19944 9904 19972
rect 8389 19935 8447 19941
rect 8404 19904 8432 19935
rect 6472 19876 8432 19904
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19805 6239 19839
rect 6181 19799 6239 19805
rect 6365 19839 6423 19845
rect 6365 19805 6377 19839
rect 6411 19805 6423 19839
rect 6365 19799 6423 19805
rect 3988 19740 4108 19768
rect 4157 19771 4215 19777
rect 3988 19712 4016 19740
rect 4157 19737 4169 19771
rect 4203 19737 4215 19771
rect 4157 19731 4215 19737
rect 4295 19771 4353 19777
rect 4295 19737 4307 19771
rect 4341 19768 4353 19771
rect 4614 19768 4620 19780
rect 4341 19740 4620 19768
rect 4341 19737 4353 19740
rect 4295 19731 4353 19737
rect 1762 19660 1768 19712
rect 1820 19660 1826 19712
rect 2958 19660 2964 19712
rect 3016 19660 3022 19712
rect 3970 19660 3976 19712
rect 4028 19660 4034 19712
rect 4172 19700 4200 19731
rect 4614 19728 4620 19740
rect 4672 19768 4678 19780
rect 6196 19768 6224 19799
rect 4672 19740 6224 19768
rect 4672 19728 4678 19740
rect 5074 19700 5080 19712
rect 4172 19672 5080 19700
rect 5074 19660 5080 19672
rect 5132 19660 5138 19712
rect 5166 19660 5172 19712
rect 5224 19660 5230 19712
rect 5629 19703 5687 19709
rect 5629 19669 5641 19703
rect 5675 19700 5687 19703
rect 5997 19703 6055 19709
rect 5997 19700 6009 19703
rect 5675 19672 6009 19700
rect 5675 19669 5687 19672
rect 5629 19663 5687 19669
rect 5997 19669 6009 19672
rect 6043 19669 6055 19703
rect 6196 19700 6224 19740
rect 6273 19771 6331 19777
rect 6273 19737 6285 19771
rect 6319 19768 6331 19771
rect 6472 19768 6500 19876
rect 8404 19848 8432 19876
rect 8496 19876 9720 19904
rect 6546 19796 6552 19848
rect 6604 19796 6610 19848
rect 6638 19796 6644 19848
rect 6696 19796 6702 19848
rect 8386 19796 8392 19848
rect 8444 19796 8450 19848
rect 6319 19740 6500 19768
rect 6319 19737 6331 19740
rect 6273 19731 6331 19737
rect 6914 19728 6920 19780
rect 6972 19728 6978 19780
rect 8294 19768 8300 19780
rect 8142 19740 8300 19768
rect 8294 19728 8300 19740
rect 8352 19728 8358 19780
rect 7558 19700 7564 19712
rect 6196 19672 7564 19700
rect 5997 19663 6055 19669
rect 7558 19660 7564 19672
rect 7616 19700 7622 19712
rect 8496 19700 8524 19876
rect 9692 19848 9720 19876
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19836 9275 19839
rect 9306 19836 9312 19848
rect 9263 19808 9312 19836
rect 9263 19805 9275 19808
rect 9217 19799 9275 19805
rect 9306 19796 9312 19808
rect 9364 19796 9370 19848
rect 9490 19796 9496 19848
rect 9548 19796 9554 19848
rect 9582 19796 9588 19848
rect 9640 19796 9646 19848
rect 9674 19796 9680 19848
rect 9732 19796 9738 19848
rect 9876 19845 9904 19944
rect 10413 19941 10425 19975
rect 10459 19972 10471 19975
rect 11790 19972 11796 19984
rect 10459 19944 11796 19972
rect 10459 19941 10471 19944
rect 10413 19935 10471 19941
rect 11790 19932 11796 19944
rect 11848 19932 11854 19984
rect 12894 19932 12900 19984
rect 12952 19972 12958 19984
rect 13446 19972 13452 19984
rect 12952 19944 13452 19972
rect 12952 19932 12958 19944
rect 13446 19932 13452 19944
rect 13504 19932 13510 19984
rect 14366 19932 14372 19984
rect 14424 19972 14430 19984
rect 15580 19972 15608 20003
rect 16114 20000 16120 20012
rect 16172 20000 16178 20052
rect 16393 20043 16451 20049
rect 16393 20009 16405 20043
rect 16439 20009 16451 20043
rect 16393 20003 16451 20009
rect 14424 19944 15608 19972
rect 14424 19932 14430 19944
rect 14752 19916 14780 19944
rect 15838 19932 15844 19984
rect 15896 19932 15902 19984
rect 16408 19972 16436 20003
rect 16850 20000 16856 20052
rect 16908 20000 16914 20052
rect 17678 20000 17684 20052
rect 17736 20000 17742 20052
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 18230 20040 18236 20052
rect 18012 20012 18236 20040
rect 18012 20000 18018 20012
rect 18230 20000 18236 20012
rect 18288 20000 18294 20052
rect 18690 20000 18696 20052
rect 18748 20040 18754 20052
rect 18877 20043 18935 20049
rect 18877 20040 18889 20043
rect 18748 20012 18889 20040
rect 18748 20000 18754 20012
rect 18877 20009 18889 20012
rect 18923 20009 18935 20043
rect 18877 20003 18935 20009
rect 20165 20043 20223 20049
rect 20165 20009 20177 20043
rect 20211 20040 20223 20043
rect 20806 20040 20812 20052
rect 20211 20012 20812 20040
rect 20211 20009 20223 20012
rect 20165 20003 20223 20009
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 22186 20000 22192 20052
rect 22244 20040 22250 20052
rect 22922 20040 22928 20052
rect 22244 20012 22928 20040
rect 22244 20000 22250 20012
rect 22922 20000 22928 20012
rect 22980 20000 22986 20052
rect 23109 20043 23167 20049
rect 23109 20009 23121 20043
rect 23155 20040 23167 20043
rect 23382 20040 23388 20052
rect 23155 20012 23388 20040
rect 23155 20009 23167 20012
rect 23109 20003 23167 20009
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 23937 20043 23995 20049
rect 23937 20009 23949 20043
rect 23983 20040 23995 20043
rect 24118 20040 24124 20052
rect 23983 20012 24124 20040
rect 23983 20009 23995 20012
rect 23937 20003 23995 20009
rect 24118 20000 24124 20012
rect 24176 20000 24182 20052
rect 26326 20000 26332 20052
rect 26384 20000 26390 20052
rect 26418 20000 26424 20052
rect 26476 20000 26482 20052
rect 28626 20000 28632 20052
rect 28684 20000 28690 20052
rect 28810 20000 28816 20052
rect 28868 20000 28874 20052
rect 28902 20000 28908 20052
rect 28960 20040 28966 20052
rect 29730 20040 29736 20052
rect 28960 20012 29736 20040
rect 28960 20000 28966 20012
rect 29730 20000 29736 20012
rect 29788 20040 29794 20052
rect 29788 20012 30052 20040
rect 29788 20000 29794 20012
rect 16574 19972 16580 19984
rect 16408 19944 16580 19972
rect 16574 19932 16580 19944
rect 16632 19932 16638 19984
rect 16669 19975 16727 19981
rect 16669 19941 16681 19975
rect 16715 19972 16727 19975
rect 17696 19972 17724 20000
rect 16715 19944 17724 19972
rect 16715 19941 16727 19944
rect 16669 19935 16727 19941
rect 17770 19932 17776 19984
rect 17828 19972 17834 19984
rect 25593 19975 25651 19981
rect 17828 19944 24164 19972
rect 17828 19932 17834 19944
rect 12161 19907 12219 19913
rect 9968 19876 10272 19904
rect 9968 19848 9996 19876
rect 9861 19839 9919 19845
rect 9861 19805 9873 19839
rect 9907 19805 9919 19839
rect 9861 19799 9919 19805
rect 9950 19796 9956 19848
rect 10008 19796 10014 19848
rect 10134 19796 10140 19848
rect 10192 19796 10198 19848
rect 10244 19845 10272 19876
rect 12161 19873 12173 19907
rect 12207 19904 12219 19907
rect 12207 19876 14688 19904
rect 12207 19873 12219 19876
rect 12161 19867 12219 19873
rect 10229 19839 10287 19845
rect 10229 19805 10241 19839
rect 10275 19805 10287 19839
rect 10229 19799 10287 19805
rect 11977 19839 12035 19845
rect 11977 19805 11989 19839
rect 12023 19836 12035 19839
rect 12066 19836 12072 19848
rect 12023 19808 12072 19836
rect 12023 19805 12035 19808
rect 11977 19799 12035 19805
rect 12066 19796 12072 19808
rect 12124 19796 12130 19848
rect 9401 19771 9459 19777
rect 9401 19737 9413 19771
rect 9447 19737 9459 19771
rect 9600 19768 9628 19796
rect 9968 19768 9996 19796
rect 9600 19740 9996 19768
rect 10045 19771 10103 19777
rect 9401 19731 9459 19737
rect 10045 19737 10057 19771
rect 10091 19737 10103 19771
rect 10045 19731 10103 19737
rect 11609 19771 11667 19777
rect 11609 19737 11621 19771
rect 11655 19768 11667 19771
rect 12176 19768 12204 19867
rect 12253 19839 12311 19845
rect 12253 19805 12265 19839
rect 12299 19836 12311 19839
rect 12526 19836 12532 19848
rect 12299 19808 12532 19836
rect 12299 19805 12311 19808
rect 12253 19799 12311 19805
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 13173 19839 13231 19845
rect 13173 19805 13185 19839
rect 13219 19836 13231 19839
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 13219 19808 13553 19836
rect 13219 19805 13231 19808
rect 13173 19799 13231 19805
rect 13541 19805 13553 19808
rect 13587 19836 13599 19839
rect 13722 19836 13728 19848
rect 13587 19808 13728 19836
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 13722 19796 13728 19808
rect 13780 19796 13786 19848
rect 13998 19796 14004 19848
rect 14056 19836 14062 19848
rect 14093 19839 14151 19845
rect 14093 19836 14105 19839
rect 14056 19808 14105 19836
rect 14056 19796 14062 19808
rect 14093 19805 14105 19808
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 14553 19839 14611 19845
rect 14553 19805 14565 19839
rect 14599 19805 14611 19839
rect 14553 19799 14611 19805
rect 11655 19740 12204 19768
rect 13265 19771 13323 19777
rect 11655 19737 11667 19740
rect 11609 19731 11667 19737
rect 13265 19737 13277 19771
rect 13311 19768 13323 19771
rect 13311 19740 13584 19768
rect 13311 19737 13323 19740
rect 13265 19731 13323 19737
rect 7616 19672 8524 19700
rect 7616 19660 7622 19672
rect 8938 19660 8944 19712
rect 8996 19700 9002 19712
rect 9416 19700 9444 19731
rect 9766 19700 9772 19712
rect 8996 19672 9772 19700
rect 8996 19660 9002 19672
rect 9766 19660 9772 19672
rect 9824 19700 9830 19712
rect 10060 19700 10088 19731
rect 9824 19672 10088 19700
rect 9824 19660 9830 19672
rect 11422 19660 11428 19712
rect 11480 19660 11486 19712
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 12713 19703 12771 19709
rect 12713 19700 12725 19703
rect 11848 19672 12725 19700
rect 11848 19660 11854 19672
rect 12713 19669 12725 19672
rect 12759 19700 12771 19703
rect 13354 19700 13360 19712
rect 12759 19672 13360 19700
rect 12759 19669 12771 19672
rect 12713 19663 12771 19669
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 13446 19660 13452 19712
rect 13504 19660 13510 19712
rect 13556 19700 13584 19740
rect 13630 19728 13636 19780
rect 13688 19768 13694 19780
rect 14568 19768 14596 19799
rect 13688 19740 14596 19768
rect 14660 19768 14688 19876
rect 14734 19864 14740 19916
rect 14792 19864 14798 19916
rect 19521 19907 19579 19913
rect 14844 19876 16988 19904
rect 14844 19768 14872 19876
rect 15197 19839 15255 19845
rect 15197 19805 15209 19839
rect 15243 19805 15255 19839
rect 15197 19799 15255 19805
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19836 15347 19839
rect 15470 19836 15476 19848
rect 15335 19808 15476 19836
rect 15335 19805 15347 19808
rect 15289 19799 15347 19805
rect 14660 19740 14872 19768
rect 15212 19768 15240 19799
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 15654 19796 15660 19848
rect 15712 19836 15718 19848
rect 16206 19836 16212 19848
rect 15712 19808 16212 19836
rect 15712 19796 15718 19808
rect 16206 19796 16212 19808
rect 16264 19796 16270 19848
rect 16298 19796 16304 19848
rect 16356 19796 16362 19848
rect 16390 19796 16396 19848
rect 16448 19796 16454 19848
rect 16850 19836 16856 19848
rect 16500 19808 16856 19836
rect 16500 19768 16528 19808
rect 16850 19796 16856 19808
rect 16908 19796 16914 19848
rect 16960 19845 16988 19876
rect 19521 19873 19533 19907
rect 19567 19904 19579 19907
rect 20070 19904 20076 19916
rect 19567 19876 20076 19904
rect 19567 19873 19579 19876
rect 19521 19867 19579 19873
rect 20070 19864 20076 19876
rect 20128 19904 20134 19916
rect 20257 19907 20315 19913
rect 20257 19904 20269 19907
rect 20128 19876 20269 19904
rect 20128 19864 20134 19876
rect 20257 19873 20269 19876
rect 20303 19873 20315 19907
rect 20257 19867 20315 19873
rect 20990 19864 20996 19916
rect 21048 19904 21054 19916
rect 23017 19907 23075 19913
rect 23017 19904 23029 19907
rect 21048 19876 23029 19904
rect 21048 19864 21054 19876
rect 23017 19873 23029 19876
rect 23063 19904 23075 19907
rect 23063 19876 23428 19904
rect 23063 19873 23075 19876
rect 23017 19867 23075 19873
rect 23400 19848 23428 19876
rect 23842 19864 23848 19916
rect 23900 19864 23906 19916
rect 23934 19864 23940 19916
rect 23992 19864 23998 19916
rect 24136 19913 24164 19944
rect 25593 19941 25605 19975
rect 25639 19972 25651 19975
rect 28644 19972 28672 20000
rect 25639 19944 28672 19972
rect 25639 19941 25651 19944
rect 25593 19935 25651 19941
rect 24121 19907 24179 19913
rect 24121 19873 24133 19907
rect 24167 19873 24179 19907
rect 24857 19907 24915 19913
rect 24857 19904 24869 19907
rect 24121 19867 24179 19873
rect 24228 19876 24869 19904
rect 16945 19839 17003 19845
rect 16945 19805 16957 19839
rect 16991 19805 17003 19839
rect 16945 19799 17003 19805
rect 17402 19796 17408 19848
rect 17460 19796 17466 19848
rect 17862 19796 17868 19848
rect 17920 19796 17926 19848
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19805 18199 19839
rect 18141 19799 18199 19805
rect 15212 19740 16528 19768
rect 13688 19728 13694 19740
rect 16574 19728 16580 19780
rect 16632 19768 16638 19780
rect 17420 19768 17448 19796
rect 16632 19740 17448 19768
rect 16632 19728 16638 19740
rect 18156 19712 18184 19799
rect 18690 19796 18696 19848
rect 18748 19796 18754 19848
rect 18961 19839 19019 19845
rect 18961 19805 18973 19839
rect 19007 19836 19019 19839
rect 19058 19836 19064 19848
rect 19007 19808 19064 19836
rect 19007 19805 19019 19808
rect 18961 19799 19019 19805
rect 19058 19796 19064 19808
rect 19116 19836 19122 19848
rect 19116 19808 19288 19836
rect 19116 19796 19122 19808
rect 19260 19780 19288 19808
rect 19886 19796 19892 19848
rect 19944 19796 19950 19848
rect 19978 19796 19984 19848
rect 20036 19796 20042 19848
rect 20346 19836 20352 19848
rect 20088 19808 20352 19836
rect 18230 19728 18236 19780
rect 18288 19728 18294 19780
rect 19242 19728 19248 19780
rect 19300 19768 19306 19780
rect 19613 19771 19671 19777
rect 19613 19768 19625 19771
rect 19300 19740 19625 19768
rect 19300 19728 19306 19740
rect 19613 19737 19625 19740
rect 19659 19768 19671 19771
rect 20088 19768 20116 19808
rect 20346 19796 20352 19808
rect 20404 19796 20410 19848
rect 20530 19796 20536 19848
rect 20588 19796 20594 19848
rect 20625 19839 20683 19845
rect 20625 19805 20637 19839
rect 20671 19805 20683 19839
rect 20625 19799 20683 19805
rect 20717 19839 20775 19845
rect 20717 19805 20729 19839
rect 20763 19836 20775 19839
rect 20901 19839 20959 19845
rect 20763 19808 20852 19836
rect 20763 19805 20775 19808
rect 20717 19799 20775 19805
rect 20640 19768 20668 19799
rect 20824 19780 20852 19808
rect 20901 19805 20913 19839
rect 20947 19805 20959 19839
rect 20901 19799 20959 19805
rect 19659 19740 20116 19768
rect 20180 19740 20668 19768
rect 19659 19737 19671 19740
rect 19613 19731 19671 19737
rect 13998 19700 14004 19712
rect 13556 19672 14004 19700
rect 13998 19660 14004 19672
rect 14056 19700 14062 19712
rect 17954 19700 17960 19712
rect 14056 19672 17960 19700
rect 14056 19660 14062 19672
rect 17954 19660 17960 19672
rect 18012 19660 18018 19712
rect 18138 19660 18144 19712
rect 18196 19660 18202 19712
rect 18248 19700 18276 19728
rect 20180 19712 20208 19740
rect 20806 19728 20812 19780
rect 20864 19728 20870 19780
rect 18874 19700 18880 19712
rect 18248 19672 18880 19700
rect 18874 19660 18880 19672
rect 18932 19660 18938 19712
rect 20162 19660 20168 19712
rect 20220 19660 20226 19712
rect 20622 19660 20628 19712
rect 20680 19700 20686 19712
rect 20916 19700 20944 19799
rect 22646 19796 22652 19848
rect 22704 19836 22710 19848
rect 23109 19839 23167 19845
rect 23109 19836 23121 19839
rect 22704 19808 23121 19836
rect 22704 19796 22710 19808
rect 23109 19805 23121 19808
rect 23155 19836 23167 19839
rect 23290 19836 23296 19848
rect 23155 19808 23296 19836
rect 23155 19805 23167 19808
rect 23109 19799 23167 19805
rect 23290 19796 23296 19808
rect 23348 19796 23354 19848
rect 23382 19796 23388 19848
rect 23440 19796 23446 19848
rect 23566 19796 23572 19848
rect 23624 19836 23630 19848
rect 23661 19839 23719 19845
rect 23661 19836 23673 19839
rect 23624 19808 23673 19836
rect 23624 19796 23630 19808
rect 23661 19805 23673 19808
rect 23707 19836 23719 19839
rect 23952 19836 23980 19864
rect 24228 19845 24256 19876
rect 24857 19873 24869 19876
rect 24903 19904 24915 19907
rect 25685 19907 25743 19913
rect 25685 19904 25697 19907
rect 24903 19876 25697 19904
rect 24903 19873 24915 19876
rect 24857 19867 24915 19873
rect 25685 19873 25697 19876
rect 25731 19873 25743 19907
rect 25685 19867 25743 19873
rect 26326 19864 26332 19916
rect 26384 19904 26390 19916
rect 28718 19904 28724 19916
rect 26384 19876 26648 19904
rect 26384 19864 26390 19876
rect 23707 19808 23980 19836
rect 24029 19839 24087 19845
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 24029 19805 24041 19839
rect 24075 19805 24087 19839
rect 24029 19799 24087 19805
rect 24213 19839 24271 19845
rect 24213 19805 24225 19839
rect 24259 19805 24271 19839
rect 24213 19799 24271 19805
rect 24397 19839 24455 19845
rect 24397 19805 24409 19839
rect 24443 19836 24455 19839
rect 24486 19836 24492 19848
rect 24443 19808 24492 19836
rect 24443 19805 24455 19808
rect 24397 19799 24455 19805
rect 22830 19728 22836 19780
rect 22888 19728 22894 19780
rect 23937 19771 23995 19777
rect 23937 19768 23949 19771
rect 23308 19740 23949 19768
rect 23308 19709 23336 19740
rect 23937 19737 23949 19740
rect 23983 19737 23995 19771
rect 23937 19731 23995 19737
rect 20680 19672 20944 19700
rect 23293 19703 23351 19709
rect 20680 19660 20686 19672
rect 23293 19669 23305 19703
rect 23339 19669 23351 19703
rect 23293 19663 23351 19669
rect 23474 19660 23480 19712
rect 23532 19660 23538 19712
rect 23566 19660 23572 19712
rect 23624 19700 23630 19712
rect 24044 19700 24072 19799
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 24581 19839 24639 19845
rect 24581 19805 24593 19839
rect 24627 19836 24639 19839
rect 24670 19836 24676 19848
rect 24627 19808 24676 19836
rect 24627 19805 24639 19808
rect 24581 19799 24639 19805
rect 24397 19703 24455 19709
rect 24397 19700 24409 19703
rect 23624 19672 24409 19700
rect 23624 19660 23630 19672
rect 24397 19669 24409 19672
rect 24443 19669 24455 19703
rect 24596 19700 24624 19799
rect 24670 19796 24676 19808
rect 24728 19796 24734 19848
rect 24762 19796 24768 19848
rect 24820 19796 24826 19848
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 25041 19839 25099 19845
rect 25041 19805 25053 19839
rect 25087 19836 25099 19839
rect 25130 19836 25136 19848
rect 25087 19808 25136 19836
rect 25087 19805 25099 19808
rect 25041 19799 25099 19805
rect 24854 19728 24860 19780
rect 24912 19768 24918 19780
rect 24964 19768 24992 19799
rect 25130 19796 25136 19808
rect 25188 19796 25194 19848
rect 25409 19839 25467 19845
rect 25409 19805 25421 19839
rect 25455 19836 25467 19839
rect 25498 19836 25504 19848
rect 25455 19808 25504 19836
rect 25455 19805 25467 19808
rect 25409 19799 25467 19805
rect 25498 19796 25504 19808
rect 25556 19796 25562 19848
rect 25866 19796 25872 19848
rect 25924 19836 25930 19848
rect 26620 19845 26648 19876
rect 28460 19876 28724 19904
rect 26053 19839 26111 19845
rect 26053 19836 26065 19839
rect 25924 19808 26065 19836
rect 25924 19796 25930 19808
rect 26053 19805 26065 19808
rect 26099 19805 26111 19839
rect 26053 19799 26111 19805
rect 26145 19839 26203 19845
rect 26145 19805 26157 19839
rect 26191 19836 26203 19839
rect 26605 19839 26663 19845
rect 26191 19808 26556 19836
rect 26191 19805 26203 19808
rect 26145 19799 26203 19805
rect 24912 19740 24992 19768
rect 24912 19728 24918 19740
rect 25222 19728 25228 19780
rect 25280 19728 25286 19780
rect 25314 19728 25320 19780
rect 25372 19728 25378 19780
rect 26528 19700 26556 19808
rect 26605 19805 26617 19839
rect 26651 19805 26663 19839
rect 26605 19799 26663 19805
rect 26694 19796 26700 19848
rect 26752 19796 26758 19848
rect 26973 19839 27031 19845
rect 26973 19805 26985 19839
rect 27019 19836 27031 19839
rect 27154 19836 27160 19848
rect 27019 19808 27160 19836
rect 27019 19805 27031 19808
rect 26973 19799 27031 19805
rect 27154 19796 27160 19808
rect 27212 19796 27218 19848
rect 27246 19796 27252 19848
rect 27304 19796 27310 19848
rect 28460 19845 28488 19876
rect 28718 19864 28724 19876
rect 28776 19864 28782 19916
rect 28445 19839 28503 19845
rect 28445 19805 28457 19839
rect 28491 19805 28503 19839
rect 28445 19799 28503 19805
rect 28629 19839 28687 19845
rect 28629 19805 28641 19839
rect 28675 19805 28687 19839
rect 28828 19836 28856 20000
rect 29089 19975 29147 19981
rect 29089 19941 29101 19975
rect 29135 19972 29147 19975
rect 29135 19944 29868 19972
rect 29135 19941 29147 19944
rect 29089 19935 29147 19941
rect 29546 19864 29552 19916
rect 29604 19864 29610 19916
rect 28905 19839 28963 19845
rect 28905 19836 28917 19839
rect 28828 19808 28917 19836
rect 28629 19799 28687 19805
rect 28905 19805 28917 19808
rect 28951 19805 28963 19839
rect 28905 19799 28963 19805
rect 29003 19839 29061 19845
rect 29003 19805 29015 19839
rect 29049 19836 29061 19839
rect 29181 19839 29239 19845
rect 29049 19808 29132 19836
rect 29049 19805 29061 19808
rect 29003 19799 29061 19805
rect 26786 19728 26792 19780
rect 26844 19728 26850 19780
rect 27264 19768 27292 19796
rect 28460 19768 28488 19799
rect 27264 19740 28488 19768
rect 28534 19728 28540 19780
rect 28592 19728 28598 19780
rect 28644 19768 28672 19799
rect 28813 19771 28871 19777
rect 28813 19768 28825 19771
rect 28644 19740 28825 19768
rect 28813 19737 28825 19740
rect 28859 19737 28871 19771
rect 29104 19768 29132 19808
rect 29181 19805 29193 19839
rect 29227 19836 29239 19839
rect 29564 19836 29592 19864
rect 29840 19848 29868 19944
rect 29227 19808 29592 19836
rect 29227 19805 29239 19808
rect 29181 19799 29239 19805
rect 29638 19796 29644 19848
rect 29696 19836 29702 19848
rect 29733 19839 29791 19845
rect 29733 19836 29745 19839
rect 29696 19808 29745 19836
rect 29696 19796 29702 19808
rect 29733 19805 29745 19808
rect 29779 19805 29791 19839
rect 29733 19799 29791 19805
rect 29822 19796 29828 19848
rect 29880 19796 29886 19848
rect 30024 19845 30052 20012
rect 30650 20000 30656 20052
rect 30708 20000 30714 20052
rect 32030 20000 32036 20052
rect 32088 20000 32094 20052
rect 34698 20000 34704 20052
rect 34756 20040 34762 20052
rect 34885 20043 34943 20049
rect 34885 20040 34897 20043
rect 34756 20012 34897 20040
rect 34756 20000 34762 20012
rect 34885 20009 34897 20012
rect 34931 20009 34943 20043
rect 34885 20003 34943 20009
rect 35158 20000 35164 20052
rect 35216 20040 35222 20052
rect 35710 20040 35716 20052
rect 35216 20012 35716 20040
rect 35216 20000 35222 20012
rect 35710 20000 35716 20012
rect 35768 20000 35774 20052
rect 35802 20000 35808 20052
rect 35860 20040 35866 20052
rect 36725 20043 36783 20049
rect 36725 20040 36737 20043
rect 35860 20012 36737 20040
rect 35860 20000 35866 20012
rect 36725 20009 36737 20012
rect 36771 20009 36783 20043
rect 36725 20003 36783 20009
rect 30116 19876 30604 19904
rect 30116 19845 30144 19876
rect 30009 19839 30067 19845
rect 30009 19805 30021 19839
rect 30055 19805 30067 19839
rect 30009 19799 30067 19805
rect 30101 19839 30159 19845
rect 30101 19805 30113 19839
rect 30147 19805 30159 19839
rect 30101 19799 30159 19805
rect 30377 19839 30435 19845
rect 30377 19805 30389 19839
rect 30423 19805 30435 19839
rect 30377 19799 30435 19805
rect 29104 19740 29224 19768
rect 28813 19731 28871 19737
rect 29196 19712 29224 19740
rect 29362 19728 29368 19780
rect 29420 19768 29426 19780
rect 30190 19768 30196 19780
rect 29420 19740 30196 19768
rect 29420 19728 29426 19740
rect 30190 19728 30196 19740
rect 30248 19768 30254 19780
rect 30392 19768 30420 19799
rect 30248 19740 30420 19768
rect 30576 19768 30604 19876
rect 30668 19845 30696 20000
rect 31036 19944 31984 19972
rect 30742 19864 30748 19916
rect 30800 19904 30806 19916
rect 31036 19913 31064 19944
rect 31021 19907 31079 19913
rect 31021 19904 31033 19907
rect 30800 19876 31033 19904
rect 30800 19864 30806 19876
rect 31021 19873 31033 19876
rect 31067 19873 31079 19907
rect 31021 19867 31079 19873
rect 31202 19864 31208 19916
rect 31260 19864 31266 19916
rect 30653 19839 30711 19845
rect 30653 19805 30665 19839
rect 30699 19805 30711 19839
rect 30653 19799 30711 19805
rect 31481 19839 31539 19845
rect 31481 19805 31493 19839
rect 31527 19836 31539 19839
rect 31570 19836 31576 19848
rect 31527 19808 31576 19836
rect 31527 19805 31539 19808
rect 31481 19799 31539 19805
rect 31496 19768 31524 19799
rect 31570 19796 31576 19808
rect 31628 19796 31634 19848
rect 31956 19845 31984 19944
rect 32048 19913 32076 20000
rect 32309 19975 32367 19981
rect 32309 19941 32321 19975
rect 32355 19972 32367 19975
rect 34606 19972 34612 19984
rect 32355 19944 34612 19972
rect 32355 19941 32367 19944
rect 32309 19935 32367 19941
rect 34606 19932 34612 19944
rect 34664 19932 34670 19984
rect 35529 19975 35587 19981
rect 35529 19941 35541 19975
rect 35575 19941 35587 19975
rect 35728 19972 35756 20000
rect 35728 19944 36584 19972
rect 35529 19935 35587 19941
rect 32033 19907 32091 19913
rect 32033 19873 32045 19907
rect 32079 19873 32091 19907
rect 32033 19867 32091 19873
rect 32950 19864 32956 19916
rect 33008 19864 33014 19916
rect 33134 19864 33140 19916
rect 33192 19904 33198 19916
rect 35544 19904 35572 19935
rect 33192 19876 33640 19904
rect 33192 19864 33198 19876
rect 31941 19839 31999 19845
rect 31941 19805 31953 19839
rect 31987 19805 31999 19839
rect 32968 19836 32996 19864
rect 33612 19845 33640 19876
rect 35084 19876 35572 19904
rect 35084 19845 35112 19876
rect 33413 19839 33471 19845
rect 33413 19836 33425 19839
rect 32968 19808 33425 19836
rect 31941 19799 31999 19805
rect 33413 19805 33425 19808
rect 33459 19805 33471 19839
rect 33413 19799 33471 19805
rect 33597 19839 33655 19845
rect 33597 19805 33609 19839
rect 33643 19805 33655 19839
rect 33597 19799 33655 19805
rect 35069 19839 35127 19845
rect 35069 19805 35081 19839
rect 35115 19805 35127 19839
rect 35069 19799 35127 19805
rect 35158 19796 35164 19848
rect 35216 19796 35222 19848
rect 35345 19839 35403 19845
rect 35345 19805 35357 19839
rect 35391 19805 35403 19839
rect 35345 19799 35403 19805
rect 30576 19740 31524 19768
rect 35360 19768 35388 19799
rect 35434 19796 35440 19848
rect 35492 19796 35498 19848
rect 35544 19836 35572 19876
rect 35618 19864 35624 19916
rect 35676 19904 35682 19916
rect 36081 19907 36139 19913
rect 36081 19904 36093 19907
rect 35676 19876 36093 19904
rect 35676 19864 35682 19876
rect 36081 19873 36093 19876
rect 36127 19873 36139 19907
rect 36081 19867 36139 19873
rect 36556 19845 36584 19944
rect 36357 19839 36415 19845
rect 36357 19836 36369 19839
rect 35544 19808 36369 19836
rect 36357 19805 36369 19808
rect 36403 19805 36415 19839
rect 36357 19799 36415 19805
rect 36541 19839 36599 19845
rect 36541 19805 36553 19839
rect 36587 19836 36599 19839
rect 36633 19839 36691 19845
rect 36633 19836 36645 19839
rect 36587 19808 36645 19836
rect 36587 19805 36599 19808
rect 36541 19799 36599 19805
rect 36633 19805 36645 19808
rect 36679 19805 36691 19839
rect 36633 19799 36691 19805
rect 36449 19771 36507 19777
rect 36449 19768 36461 19771
rect 35360 19740 36461 19768
rect 30248 19728 30254 19740
rect 36449 19737 36461 19740
rect 36495 19737 36507 19771
rect 36449 19731 36507 19737
rect 28948 19700 28954 19712
rect 24596 19672 28954 19700
rect 24397 19663 24455 19669
rect 28948 19660 28954 19672
rect 29006 19660 29012 19712
rect 29178 19660 29184 19712
rect 29236 19660 29242 19712
rect 29546 19660 29552 19712
rect 29604 19660 29610 19712
rect 33505 19703 33563 19709
rect 33505 19669 33517 19703
rect 33551 19700 33563 19703
rect 34790 19700 34796 19712
rect 33551 19672 34796 19700
rect 33551 19669 33563 19672
rect 33505 19663 33563 19669
rect 34790 19660 34796 19672
rect 34848 19660 34854 19712
rect 35894 19660 35900 19712
rect 35952 19660 35958 19712
rect 35989 19703 36047 19709
rect 35989 19669 36001 19703
rect 36035 19700 36047 19703
rect 36170 19700 36176 19712
rect 36035 19672 36176 19700
rect 36035 19669 36047 19672
rect 35989 19663 36047 19669
rect 36170 19660 36176 19672
rect 36228 19660 36234 19712
rect 1104 19610 38272 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38272 19610
rect 1104 19536 38272 19558
rect 1394 19456 1400 19508
rect 1452 19496 1458 19508
rect 1452 19468 4016 19496
rect 1452 19456 1458 19468
rect 1412 19369 1440 19456
rect 1673 19431 1731 19437
rect 1673 19397 1685 19431
rect 1719 19428 1731 19431
rect 1762 19428 1768 19440
rect 1719 19400 1768 19428
rect 1719 19397 1731 19400
rect 1673 19391 1731 19397
rect 1762 19388 1768 19400
rect 1820 19388 1826 19440
rect 2958 19428 2964 19440
rect 2898 19400 2964 19428
rect 2958 19388 2964 19400
rect 3016 19428 3022 19440
rect 3016 19400 3832 19428
rect 3016 19388 3022 19400
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19329 1455 19363
rect 1397 19323 1455 19329
rect 3513 19363 3571 19369
rect 3513 19329 3525 19363
rect 3559 19360 3571 19363
rect 3602 19360 3608 19372
rect 3559 19332 3608 19360
rect 3559 19329 3571 19332
rect 3513 19323 3571 19329
rect 3602 19320 3608 19332
rect 3660 19320 3666 19372
rect 3697 19363 3755 19369
rect 3697 19329 3709 19363
rect 3743 19329 3755 19363
rect 3804 19360 3832 19400
rect 3878 19388 3884 19440
rect 3936 19388 3942 19440
rect 3988 19360 4016 19468
rect 5074 19456 5080 19508
rect 5132 19496 5138 19508
rect 5132 19468 5764 19496
rect 5132 19456 5138 19468
rect 5736 19428 5764 19468
rect 5902 19456 5908 19508
rect 5960 19456 5966 19508
rect 6546 19456 6552 19508
rect 6604 19456 6610 19508
rect 6914 19456 6920 19508
rect 6972 19496 6978 19508
rect 7009 19499 7067 19505
rect 7009 19496 7021 19499
rect 6972 19468 7021 19496
rect 6972 19456 6978 19468
rect 7009 19465 7021 19468
rect 7055 19465 7067 19499
rect 7009 19459 7067 19465
rect 7190 19456 7196 19508
rect 7248 19456 7254 19508
rect 8202 19456 8208 19508
rect 8260 19496 8266 19508
rect 9309 19499 9367 19505
rect 9309 19496 9321 19499
rect 8260 19468 9321 19496
rect 8260 19456 8266 19468
rect 9309 19465 9321 19468
rect 9355 19465 9367 19499
rect 9309 19459 9367 19465
rect 9582 19456 9588 19508
rect 9640 19456 9646 19508
rect 11790 19496 11796 19508
rect 9692 19468 11796 19496
rect 6564 19428 6592 19456
rect 5736 19400 6592 19428
rect 4157 19363 4215 19369
rect 4157 19360 4169 19363
rect 3804 19332 3924 19360
rect 3697 19323 3755 19329
rect 3712 19292 3740 19323
rect 3160 19264 3740 19292
rect 3160 19236 3188 19264
rect 3142 19184 3148 19236
rect 3200 19184 3206 19236
rect 3896 19224 3924 19332
rect 3988 19332 4169 19360
rect 3988 19304 4016 19332
rect 4157 19329 4169 19332
rect 4203 19329 4215 19363
rect 4157 19323 4215 19329
rect 5442 19320 5448 19372
rect 5500 19360 5506 19372
rect 7208 19369 7236 19456
rect 8938 19388 8944 19440
rect 8996 19388 9002 19440
rect 9030 19388 9036 19440
rect 9088 19388 9094 19440
rect 9600 19428 9628 19456
rect 9140 19400 9628 19428
rect 7193 19363 7251 19369
rect 5500 19332 7144 19360
rect 5500 19320 5506 19332
rect 3970 19252 3976 19304
rect 4028 19252 4034 19304
rect 4433 19295 4491 19301
rect 4433 19261 4445 19295
rect 4479 19292 4491 19295
rect 4798 19292 4804 19304
rect 4479 19264 4804 19292
rect 4479 19261 4491 19264
rect 4433 19255 4491 19261
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 3896 19196 4016 19224
rect 3988 19156 4016 19196
rect 5460 19156 5488 19320
rect 7116 19292 7144 19332
rect 7193 19329 7205 19363
rect 7239 19329 7251 19363
rect 7929 19363 7987 19369
rect 7929 19360 7941 19363
rect 7193 19323 7251 19329
rect 7300 19332 7941 19360
rect 7300 19292 7328 19332
rect 7929 19329 7941 19332
rect 7975 19360 7987 19363
rect 8202 19360 8208 19372
rect 7975 19332 8208 19360
rect 7975 19329 7987 19332
rect 7929 19323 7987 19329
rect 8202 19320 8208 19332
rect 8260 19320 8266 19372
rect 8754 19320 8760 19372
rect 8812 19320 8818 19372
rect 9140 19369 9168 19400
rect 9125 19363 9183 19369
rect 9125 19329 9137 19363
rect 9171 19329 9183 19363
rect 9125 19323 9183 19329
rect 9490 19320 9496 19372
rect 9548 19360 9554 19372
rect 9585 19363 9643 19369
rect 9585 19360 9597 19363
rect 9548 19332 9597 19360
rect 9548 19320 9554 19332
rect 9585 19329 9597 19332
rect 9631 19360 9643 19363
rect 9692 19360 9720 19468
rect 11790 19456 11796 19468
rect 11848 19456 11854 19508
rect 12345 19499 12403 19505
rect 12345 19496 12357 19499
rect 11992 19468 12357 19496
rect 11164 19400 11560 19428
rect 9631 19332 9720 19360
rect 9769 19363 9827 19369
rect 9631 19329 9643 19332
rect 9585 19323 9643 19329
rect 9769 19329 9781 19363
rect 9815 19360 9827 19363
rect 9950 19360 9956 19372
rect 9815 19332 9956 19360
rect 9815 19329 9827 19332
rect 9769 19323 9827 19329
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 11164 19369 11192 19400
rect 11532 19369 11560 19400
rect 11149 19363 11207 19369
rect 11149 19360 11161 19363
rect 11112 19332 11161 19360
rect 11112 19320 11118 19332
rect 11149 19329 11161 19332
rect 11195 19329 11207 19363
rect 11149 19323 11207 19329
rect 11333 19363 11391 19369
rect 11333 19329 11345 19363
rect 11379 19360 11391 19363
rect 11517 19363 11575 19369
rect 11379 19332 11413 19360
rect 11379 19329 11391 19332
rect 11333 19323 11391 19329
rect 11517 19329 11529 19363
rect 11563 19329 11575 19363
rect 11517 19323 11575 19329
rect 7116 19264 7328 19292
rect 8294 19252 8300 19304
rect 8352 19252 8358 19304
rect 9306 19252 9312 19304
rect 9364 19292 9370 19304
rect 9401 19295 9459 19301
rect 9401 19292 9413 19295
rect 9364 19264 9413 19292
rect 9364 19252 9370 19264
rect 9401 19261 9413 19264
rect 9447 19261 9459 19295
rect 11348 19292 11376 19323
rect 11882 19320 11888 19372
rect 11940 19320 11946 19372
rect 11992 19369 12020 19468
rect 12345 19465 12357 19468
rect 12391 19465 12403 19499
rect 12345 19459 12403 19465
rect 13170 19456 13176 19508
rect 13228 19456 13234 19508
rect 15654 19496 15660 19508
rect 14481 19468 15660 19496
rect 12158 19388 12164 19440
rect 12216 19428 12222 19440
rect 12989 19431 13047 19437
rect 12989 19428 13001 19431
rect 12216 19400 13001 19428
rect 12216 19388 12222 19400
rect 12989 19397 13001 19400
rect 13035 19428 13047 19431
rect 13722 19428 13728 19440
rect 13035 19400 13728 19428
rect 13035 19397 13047 19400
rect 12989 19391 13047 19397
rect 13722 19388 13728 19400
rect 13780 19388 13786 19440
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19329 12035 19363
rect 11977 19323 12035 19329
rect 12250 19320 12256 19372
rect 12308 19320 12314 19372
rect 12526 19320 12532 19372
rect 12584 19320 12590 19372
rect 12621 19363 12679 19369
rect 12621 19329 12633 19363
rect 12667 19329 12679 19363
rect 12621 19323 12679 19329
rect 11348 19264 11744 19292
rect 9401 19255 9459 19261
rect 9214 19184 9220 19236
rect 9272 19224 9278 19236
rect 11716 19233 11744 19264
rect 11790 19252 11796 19304
rect 11848 19252 11854 19304
rect 12066 19252 12072 19304
rect 12124 19292 12130 19304
rect 12636 19292 12664 19323
rect 13354 19320 13360 19372
rect 13412 19320 13418 19372
rect 14274 19320 14280 19372
rect 14332 19320 14338 19372
rect 14481 19350 14509 19468
rect 15654 19456 15660 19468
rect 15712 19456 15718 19508
rect 15838 19456 15844 19508
rect 15896 19456 15902 19508
rect 16206 19456 16212 19508
rect 16264 19496 16270 19508
rect 16264 19468 18092 19496
rect 16264 19456 16270 19468
rect 14553 19363 14611 19369
rect 14553 19350 14565 19363
rect 14481 19329 14565 19350
rect 14599 19329 14611 19363
rect 14481 19323 14611 19329
rect 14481 19322 14596 19323
rect 14734 19320 14740 19372
rect 14792 19320 14798 19372
rect 15856 19360 15884 19456
rect 16298 19388 16304 19440
rect 16356 19428 16362 19440
rect 18064 19428 18092 19468
rect 18138 19456 18144 19508
rect 18196 19496 18202 19508
rect 19518 19496 19524 19508
rect 18196 19468 19524 19496
rect 18196 19456 18202 19468
rect 19518 19456 19524 19468
rect 19576 19456 19582 19508
rect 19797 19499 19855 19505
rect 19797 19465 19809 19499
rect 19843 19496 19855 19499
rect 19978 19496 19984 19508
rect 19843 19468 19984 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 22094 19456 22100 19508
rect 22152 19496 22158 19508
rect 22649 19499 22707 19505
rect 22152 19468 22508 19496
rect 22152 19456 22158 19468
rect 19242 19428 19248 19440
rect 16356 19400 17172 19428
rect 16356 19388 16362 19400
rect 17144 19369 17172 19400
rect 17420 19400 17632 19428
rect 18064 19400 19248 19428
rect 17420 19372 17448 19400
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 15856 19332 16681 19360
rect 16669 19329 16681 19332
rect 16715 19329 16727 19363
rect 16669 19323 16727 19329
rect 17129 19363 17187 19369
rect 17129 19329 17141 19363
rect 17175 19329 17187 19363
rect 17129 19323 17187 19329
rect 17402 19320 17408 19372
rect 17460 19320 17466 19372
rect 17604 19369 17632 19400
rect 19242 19388 19248 19400
rect 19300 19388 19306 19440
rect 19536 19428 19564 19456
rect 19536 19400 19932 19428
rect 17589 19363 17647 19369
rect 17589 19329 17601 19363
rect 17635 19329 17647 19363
rect 17589 19323 17647 19329
rect 18141 19363 18199 19369
rect 18141 19329 18153 19363
rect 18187 19360 18199 19363
rect 19334 19360 19340 19372
rect 18187 19332 19340 19360
rect 18187 19329 18199 19332
rect 18141 19323 18199 19329
rect 19334 19320 19340 19332
rect 19392 19320 19398 19372
rect 19610 19320 19616 19372
rect 19668 19360 19674 19372
rect 19904 19369 19932 19400
rect 21910 19388 21916 19440
rect 21968 19428 21974 19440
rect 22189 19431 22247 19437
rect 22189 19428 22201 19431
rect 21968 19400 22201 19428
rect 21968 19388 21974 19400
rect 22189 19397 22201 19400
rect 22235 19397 22247 19431
rect 22370 19428 22376 19440
rect 22189 19391 22247 19397
rect 22296 19400 22376 19428
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19668 19332 19717 19360
rect 19668 19320 19674 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 19978 19320 19984 19372
rect 20036 19360 20042 19372
rect 20530 19360 20536 19372
rect 20036 19332 20536 19360
rect 20036 19320 20042 19332
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 12124 19264 12664 19292
rect 13541 19295 13599 19301
rect 12124 19252 12130 19264
rect 13541 19261 13553 19295
rect 13587 19292 13599 19295
rect 13906 19292 13912 19304
rect 13587 19264 13912 19292
rect 13587 19261 13599 19264
rect 13541 19255 13599 19261
rect 13906 19252 13912 19264
rect 13964 19252 13970 19304
rect 14108 19264 17080 19292
rect 11701 19227 11759 19233
rect 9272 19196 11652 19224
rect 9272 19184 9278 19196
rect 3988 19128 5488 19156
rect 11330 19116 11336 19168
rect 11388 19116 11394 19168
rect 11624 19156 11652 19196
rect 11701 19193 11713 19227
rect 11747 19224 11759 19227
rect 12158 19224 12164 19236
rect 11747 19196 12164 19224
rect 11747 19193 11759 19196
rect 11701 19187 11759 19193
rect 12158 19184 12164 19196
rect 12216 19184 12222 19236
rect 14108 19224 14136 19264
rect 12268 19196 14136 19224
rect 12268 19156 12296 19196
rect 14642 19184 14648 19236
rect 14700 19184 14706 19236
rect 16758 19184 16764 19236
rect 16816 19184 16822 19236
rect 17052 19224 17080 19264
rect 17770 19252 17776 19304
rect 17828 19292 17834 19304
rect 17957 19295 18015 19301
rect 17957 19292 17969 19295
rect 17828 19264 17969 19292
rect 17828 19252 17834 19264
rect 17957 19261 17969 19264
rect 18003 19292 18015 19295
rect 20162 19292 20168 19304
rect 18003 19264 20168 19292
rect 18003 19261 18015 19264
rect 17957 19255 18015 19261
rect 20162 19252 20168 19264
rect 20220 19252 20226 19304
rect 22296 19301 22324 19400
rect 22370 19388 22376 19400
rect 22428 19388 22434 19440
rect 22480 19369 22508 19468
rect 22649 19465 22661 19499
rect 22695 19496 22707 19499
rect 22830 19496 22836 19508
rect 22695 19468 22836 19496
rect 22695 19465 22707 19468
rect 22649 19459 22707 19465
rect 22830 19456 22836 19468
rect 22888 19456 22894 19508
rect 23842 19456 23848 19508
rect 23900 19456 23906 19508
rect 23934 19456 23940 19508
rect 23992 19496 23998 19508
rect 24762 19496 24768 19508
rect 23992 19468 24768 19496
rect 23992 19456 23998 19468
rect 24762 19456 24768 19468
rect 24820 19456 24826 19508
rect 25866 19456 25872 19508
rect 25924 19496 25930 19508
rect 27154 19496 27160 19508
rect 25924 19468 27160 19496
rect 25924 19456 25930 19468
rect 27154 19456 27160 19468
rect 27212 19456 27218 19508
rect 27801 19499 27859 19505
rect 27801 19465 27813 19499
rect 27847 19496 27859 19499
rect 28074 19496 28080 19508
rect 27847 19468 28080 19496
rect 27847 19465 27859 19468
rect 27801 19459 27859 19465
rect 28074 19456 28080 19468
rect 28132 19456 28138 19508
rect 28718 19456 28724 19508
rect 28776 19496 28782 19508
rect 29178 19496 29184 19508
rect 28776 19468 29184 19496
rect 28776 19456 28782 19468
rect 29178 19456 29184 19468
rect 29236 19456 29242 19508
rect 29546 19456 29552 19508
rect 29604 19456 29610 19508
rect 29730 19456 29736 19508
rect 29788 19456 29794 19508
rect 29822 19456 29828 19508
rect 29880 19456 29886 19508
rect 30193 19499 30251 19505
rect 30193 19465 30205 19499
rect 30239 19496 30251 19499
rect 30374 19496 30380 19508
rect 30239 19468 30380 19496
rect 30239 19465 30251 19468
rect 30193 19459 30251 19465
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 32950 19456 32956 19508
rect 33008 19496 33014 19508
rect 33781 19499 33839 19505
rect 33008 19468 33364 19496
rect 33008 19456 33014 19468
rect 23474 19388 23480 19440
rect 23532 19428 23538 19440
rect 23569 19431 23627 19437
rect 23569 19428 23581 19431
rect 23532 19400 23581 19428
rect 23532 19388 23538 19400
rect 23569 19397 23581 19400
rect 23615 19428 23627 19431
rect 24486 19428 24492 19440
rect 23615 19400 24492 19428
rect 23615 19397 23627 19400
rect 23569 19391 23627 19397
rect 22465 19363 22523 19369
rect 22465 19329 22477 19363
rect 22511 19329 22523 19363
rect 22465 19323 22523 19329
rect 22554 19320 22560 19372
rect 22612 19360 22618 19372
rect 22741 19363 22799 19369
rect 22741 19360 22753 19363
rect 22612 19332 22753 19360
rect 22612 19320 22618 19332
rect 22741 19329 22753 19332
rect 22787 19329 22799 19363
rect 22741 19323 22799 19329
rect 23106 19320 23112 19372
rect 23164 19360 23170 19372
rect 23382 19360 23388 19372
rect 23164 19332 23388 19360
rect 23164 19320 23170 19332
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 24044 19369 24072 19400
rect 24486 19388 24492 19400
rect 24544 19428 24550 19440
rect 27062 19428 27068 19440
rect 24544 19400 27068 19428
rect 24544 19388 24550 19400
rect 27062 19388 27068 19400
rect 27120 19388 27126 19440
rect 27430 19388 27436 19440
rect 27488 19388 27494 19440
rect 27522 19388 27528 19440
rect 27580 19428 27586 19440
rect 27580 19400 27625 19428
rect 27580 19388 27586 19400
rect 27982 19388 27988 19440
rect 28040 19428 28046 19440
rect 29564 19428 29592 19456
rect 28040 19400 29040 19428
rect 28040 19388 28046 19400
rect 24029 19363 24087 19369
rect 24029 19329 24041 19363
rect 24075 19360 24087 19363
rect 24075 19332 24109 19360
rect 24075 19329 24087 19332
rect 24029 19323 24087 19329
rect 27246 19320 27252 19372
rect 27304 19369 27310 19372
rect 27304 19363 27327 19369
rect 27315 19329 27327 19363
rect 27304 19323 27327 19329
rect 27304 19320 27310 19323
rect 22281 19295 22339 19301
rect 22281 19261 22293 19295
rect 22327 19261 22339 19295
rect 22281 19255 22339 19261
rect 24302 19252 24308 19304
rect 24360 19292 24366 19304
rect 27448 19292 27476 19388
rect 24360 19264 27476 19292
rect 27540 19292 27568 19388
rect 27614 19320 27620 19372
rect 27672 19320 27678 19372
rect 27798 19320 27804 19372
rect 27856 19360 27862 19372
rect 27893 19363 27951 19369
rect 27893 19360 27905 19363
rect 27856 19332 27905 19360
rect 27856 19320 27862 19332
rect 27893 19329 27905 19332
rect 27939 19329 27951 19363
rect 27893 19323 27951 19329
rect 28074 19320 28080 19372
rect 28132 19320 28138 19372
rect 28258 19320 28264 19372
rect 28316 19320 28322 19372
rect 28534 19320 28540 19372
rect 28592 19320 28598 19372
rect 29012 19369 29040 19400
rect 29196 19400 29592 19428
rect 29196 19369 29224 19400
rect 28997 19363 29055 19369
rect 28997 19329 29009 19363
rect 29043 19329 29055 19363
rect 28997 19323 29055 19329
rect 29181 19363 29239 19369
rect 29181 19329 29193 19363
rect 29227 19329 29239 19363
rect 29181 19323 29239 19329
rect 29362 19320 29368 19372
rect 29420 19320 29426 19372
rect 29457 19363 29515 19369
rect 29457 19329 29469 19363
rect 29503 19360 29515 19363
rect 29546 19360 29552 19372
rect 29503 19332 29552 19360
rect 29503 19329 29515 19332
rect 29457 19323 29515 19329
rect 29546 19320 29552 19332
rect 29604 19320 29610 19372
rect 29748 19369 29776 19456
rect 29840 19428 29868 19456
rect 29840 19400 30236 19428
rect 30208 19369 30236 19400
rect 29733 19363 29791 19369
rect 29733 19329 29745 19363
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 29825 19363 29883 19369
rect 29825 19329 29837 19363
rect 29871 19360 29883 19363
rect 30009 19363 30067 19369
rect 30009 19360 30021 19363
rect 29871 19332 30021 19360
rect 29871 19329 29883 19332
rect 29825 19323 29883 19329
rect 30009 19329 30021 19332
rect 30055 19329 30067 19363
rect 30009 19323 30067 19329
rect 30193 19363 30251 19369
rect 30193 19329 30205 19363
rect 30239 19329 30251 19363
rect 30193 19323 30251 19329
rect 32953 19363 33011 19369
rect 32953 19329 32965 19363
rect 32999 19360 33011 19363
rect 33060 19360 33088 19468
rect 33336 19437 33364 19468
rect 33781 19465 33793 19499
rect 33827 19465 33839 19499
rect 33781 19459 33839 19465
rect 33965 19499 34023 19505
rect 33965 19465 33977 19499
rect 34011 19496 34023 19499
rect 34011 19468 34560 19496
rect 34011 19465 34023 19468
rect 33965 19459 34023 19465
rect 33321 19431 33379 19437
rect 33321 19397 33333 19431
rect 33367 19397 33379 19431
rect 33796 19428 33824 19459
rect 33796 19400 34468 19428
rect 33321 19391 33379 19397
rect 32999 19332 33088 19360
rect 32999 19329 33011 19332
rect 32953 19323 33011 19329
rect 33134 19320 33140 19372
rect 33192 19320 33198 19372
rect 33873 19363 33931 19369
rect 33873 19360 33885 19363
rect 33704 19332 33885 19360
rect 28166 19292 28172 19304
rect 27540 19264 28172 19292
rect 24360 19252 24366 19264
rect 28166 19252 28172 19264
rect 28224 19252 28230 19304
rect 28552 19292 28580 19320
rect 29273 19295 29331 19301
rect 29273 19292 29285 19295
rect 28552 19264 29285 19292
rect 29273 19261 29285 19264
rect 29319 19261 29331 19295
rect 29273 19255 29331 19261
rect 25682 19224 25688 19236
rect 17052 19196 25688 19224
rect 11624 19128 12296 19156
rect 12894 19116 12900 19168
rect 12952 19116 12958 19168
rect 17218 19116 17224 19168
rect 17276 19156 17282 19168
rect 22094 19156 22100 19168
rect 17276 19128 22100 19156
rect 17276 19116 17282 19128
rect 22094 19116 22100 19128
rect 22152 19116 22158 19168
rect 22480 19165 22508 19196
rect 25682 19184 25688 19196
rect 25740 19184 25746 19236
rect 33152 19224 33180 19320
rect 33597 19227 33655 19233
rect 33597 19224 33609 19227
rect 33152 19196 33609 19224
rect 33597 19193 33609 19196
rect 33643 19193 33655 19227
rect 33597 19187 33655 19193
rect 22465 19159 22523 19165
rect 22465 19125 22477 19159
rect 22511 19125 22523 19159
rect 22465 19119 22523 19125
rect 24118 19116 24124 19168
rect 24176 19156 24182 19168
rect 24213 19159 24271 19165
rect 24213 19156 24225 19159
rect 24176 19128 24225 19156
rect 24176 19116 24182 19128
rect 24213 19125 24225 19128
rect 24259 19156 24271 19159
rect 26786 19156 26792 19168
rect 24259 19128 26792 19156
rect 24259 19125 24271 19128
rect 24213 19119 24271 19125
rect 26786 19116 26792 19128
rect 26844 19116 26850 19168
rect 29638 19116 29644 19168
rect 29696 19116 29702 19168
rect 33134 19116 33140 19168
rect 33192 19156 33198 19168
rect 33704 19156 33732 19332
rect 33873 19329 33885 19332
rect 33919 19329 33931 19363
rect 33873 19323 33931 19329
rect 34146 19320 34152 19372
rect 34204 19320 34210 19372
rect 34440 19369 34468 19400
rect 34241 19363 34299 19369
rect 34241 19329 34253 19363
rect 34287 19360 34299 19363
rect 34425 19363 34483 19369
rect 34287 19332 34376 19360
rect 34287 19329 34299 19332
rect 34241 19323 34299 19329
rect 34348 19292 34376 19332
rect 34425 19329 34437 19363
rect 34471 19329 34483 19363
rect 34532 19360 34560 19468
rect 34790 19456 34796 19508
rect 34848 19456 34854 19508
rect 35894 19456 35900 19508
rect 35952 19456 35958 19508
rect 34808 19428 34836 19456
rect 34808 19400 36032 19428
rect 34701 19363 34759 19369
rect 34701 19360 34713 19363
rect 34532 19332 34713 19360
rect 34425 19323 34483 19329
rect 34701 19329 34713 19332
rect 34747 19329 34759 19363
rect 34808 19360 34836 19400
rect 36004 19369 36032 19400
rect 34885 19363 34943 19369
rect 34885 19360 34897 19363
rect 34808 19332 34897 19360
rect 34701 19323 34759 19329
rect 34885 19329 34897 19332
rect 34931 19329 34943 19363
rect 35805 19363 35863 19369
rect 35805 19360 35817 19363
rect 34885 19323 34943 19329
rect 34992 19332 35817 19360
rect 34790 19292 34796 19304
rect 34348 19264 34796 19292
rect 34790 19252 34796 19264
rect 34848 19252 34854 19304
rect 34992 19292 35020 19332
rect 35805 19329 35817 19332
rect 35851 19329 35863 19363
rect 35805 19323 35863 19329
rect 35989 19363 36047 19369
rect 35989 19329 36001 19363
rect 36035 19329 36047 19363
rect 35989 19323 36047 19329
rect 34900 19264 35020 19292
rect 34422 19184 34428 19236
rect 34480 19224 34486 19236
rect 34900 19224 34928 19264
rect 34480 19196 34928 19224
rect 34480 19184 34486 19196
rect 33192 19128 33732 19156
rect 34609 19159 34667 19165
rect 33192 19116 33198 19128
rect 34609 19125 34621 19159
rect 34655 19156 34667 19159
rect 35986 19156 35992 19168
rect 34655 19128 35992 19156
rect 34655 19125 34667 19128
rect 34609 19119 34667 19125
rect 35986 19116 35992 19128
rect 36044 19116 36050 19168
rect 1104 19066 38272 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38272 19066
rect 1104 18992 38272 19014
rect 4709 18955 4767 18961
rect 4709 18921 4721 18955
rect 4755 18952 4767 18955
rect 4798 18952 4804 18964
rect 4755 18924 4804 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 17218 18952 17224 18964
rect 4908 18924 17224 18952
rect 4908 18884 4936 18924
rect 17218 18912 17224 18924
rect 17276 18912 17282 18964
rect 18046 18912 18052 18964
rect 18104 18952 18110 18964
rect 18966 18952 18972 18964
rect 18104 18924 18972 18952
rect 18104 18912 18110 18924
rect 18966 18912 18972 18924
rect 19024 18952 19030 18964
rect 19024 18924 19334 18952
rect 19024 18912 19030 18924
rect 13906 18884 13912 18896
rect 3160 18856 4936 18884
rect 6104 18856 13912 18884
rect 3160 18825 3188 18856
rect 3145 18819 3203 18825
rect 3145 18785 3157 18819
rect 3191 18785 3203 18819
rect 3145 18779 3203 18785
rect 3329 18819 3387 18825
rect 3329 18785 3341 18819
rect 3375 18816 3387 18819
rect 4062 18816 4068 18828
rect 3375 18788 4068 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 5721 18819 5779 18825
rect 5721 18785 5733 18819
rect 5767 18816 5779 18819
rect 5902 18816 5908 18828
rect 5767 18788 5908 18816
rect 5767 18785 5779 18788
rect 5721 18779 5779 18785
rect 5902 18776 5908 18788
rect 5960 18776 5966 18828
rect 6104 18825 6132 18856
rect 13906 18844 13912 18856
rect 13964 18884 13970 18896
rect 17865 18887 17923 18893
rect 13964 18856 14412 18884
rect 13964 18844 13970 18856
rect 6089 18819 6147 18825
rect 6089 18785 6101 18819
rect 6135 18785 6147 18819
rect 6089 18779 6147 18785
rect 10870 18776 10876 18828
rect 10928 18776 10934 18828
rect 11422 18776 11428 18828
rect 11480 18776 11486 18828
rect 11808 18788 12388 18816
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18748 4951 18751
rect 5166 18748 5172 18760
rect 4939 18720 5172 18748
rect 4939 18717 4951 18720
rect 4893 18711 4951 18717
rect 5166 18708 5172 18720
rect 5224 18708 5230 18760
rect 5994 18708 6000 18760
rect 6052 18708 6058 18760
rect 10781 18751 10839 18757
rect 10781 18717 10793 18751
rect 10827 18748 10839 18751
rect 11440 18748 11468 18776
rect 11808 18757 11836 18788
rect 12360 18760 12388 18788
rect 10827 18720 11468 18748
rect 11793 18751 11851 18757
rect 10827 18717 10839 18720
rect 10781 18711 10839 18717
rect 11793 18717 11805 18751
rect 11839 18717 11851 18751
rect 11793 18711 11851 18717
rect 11882 18708 11888 18760
rect 11940 18708 11946 18760
rect 11977 18751 12035 18757
rect 11977 18717 11989 18751
rect 12023 18748 12035 18751
rect 12066 18748 12072 18760
rect 12023 18720 12072 18748
rect 12023 18717 12035 18720
rect 11977 18711 12035 18717
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 12161 18751 12219 18757
rect 12161 18717 12173 18751
rect 12207 18717 12219 18751
rect 12161 18711 12219 18717
rect 934 18640 940 18692
rect 992 18680 998 18692
rect 1397 18683 1455 18689
rect 1397 18680 1409 18683
rect 992 18652 1409 18680
rect 992 18640 998 18652
rect 1397 18649 1409 18652
rect 1443 18649 1455 18683
rect 1397 18643 1455 18649
rect 1762 18640 1768 18692
rect 1820 18640 1826 18692
rect 3053 18683 3111 18689
rect 3053 18649 3065 18683
rect 3099 18680 3111 18683
rect 3142 18680 3148 18692
rect 3099 18652 3148 18680
rect 3099 18649 3111 18652
rect 3053 18643 3111 18649
rect 3142 18640 3148 18652
rect 3200 18640 3206 18692
rect 5626 18640 5632 18692
rect 5684 18680 5690 18692
rect 5810 18680 5816 18692
rect 5684 18652 5816 18680
rect 5684 18640 5690 18652
rect 5810 18640 5816 18652
rect 5868 18680 5874 18692
rect 9214 18680 9220 18692
rect 5868 18652 9220 18680
rect 5868 18640 5874 18652
rect 9214 18640 9220 18652
rect 9272 18640 9278 18692
rect 10689 18683 10747 18689
rect 10689 18649 10701 18683
rect 10735 18680 10747 18683
rect 11517 18683 11575 18689
rect 11517 18680 11529 18683
rect 10735 18652 11529 18680
rect 10735 18649 10747 18652
rect 10689 18643 10747 18649
rect 11517 18649 11529 18652
rect 11563 18649 11575 18683
rect 11517 18643 11575 18649
rect 1946 18572 1952 18624
rect 2004 18612 2010 18624
rect 2685 18615 2743 18621
rect 2685 18612 2697 18615
rect 2004 18584 2697 18612
rect 2004 18572 2010 18584
rect 2685 18581 2697 18584
rect 2731 18581 2743 18615
rect 2685 18575 2743 18581
rect 4246 18572 4252 18624
rect 4304 18612 4310 18624
rect 6273 18615 6331 18621
rect 6273 18612 6285 18615
rect 4304 18584 6285 18612
rect 4304 18572 4310 18584
rect 6273 18581 6285 18584
rect 6319 18581 6331 18615
rect 6273 18575 6331 18581
rect 6546 18572 6552 18624
rect 6604 18612 6610 18624
rect 6730 18612 6736 18624
rect 6604 18584 6736 18612
rect 6604 18572 6610 18584
rect 6730 18572 6736 18584
rect 6788 18612 6794 18624
rect 10042 18612 10048 18624
rect 6788 18584 10048 18612
rect 6788 18572 6794 18584
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 10318 18572 10324 18624
rect 10376 18572 10382 18624
rect 11330 18572 11336 18624
rect 11388 18612 11394 18624
rect 12176 18612 12204 18711
rect 12342 18708 12348 18760
rect 12400 18708 12406 18760
rect 14384 18757 14412 18856
rect 17865 18853 17877 18887
rect 17911 18884 17923 18887
rect 18325 18887 18383 18893
rect 18325 18884 18337 18887
rect 17911 18856 18337 18884
rect 17911 18853 17923 18856
rect 17865 18847 17923 18853
rect 18325 18853 18337 18856
rect 18371 18853 18383 18887
rect 18325 18847 18383 18853
rect 18598 18844 18604 18896
rect 18656 18844 18662 18896
rect 19306 18884 19334 18924
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 19484 18924 19809 18952
rect 19484 18912 19490 18924
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 19797 18915 19855 18921
rect 19978 18912 19984 18964
rect 20036 18912 20042 18964
rect 20162 18912 20168 18964
rect 20220 18912 20226 18964
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 20809 18955 20867 18961
rect 20809 18952 20821 18955
rect 20772 18924 20821 18952
rect 20772 18912 20778 18924
rect 20809 18921 20821 18924
rect 20855 18921 20867 18955
rect 20809 18915 20867 18921
rect 20898 18912 20904 18964
rect 20956 18952 20962 18964
rect 20993 18955 21051 18961
rect 20993 18952 21005 18955
rect 20956 18924 21005 18952
rect 20956 18912 20962 18924
rect 20993 18921 21005 18924
rect 21039 18952 21051 18955
rect 21082 18952 21088 18964
rect 21039 18924 21088 18952
rect 21039 18921 21051 18924
rect 20993 18915 21051 18921
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 22557 18955 22615 18961
rect 22557 18921 22569 18955
rect 22603 18952 22615 18955
rect 22646 18952 22652 18964
rect 22603 18924 22652 18952
rect 22603 18921 22615 18924
rect 22557 18915 22615 18921
rect 22646 18912 22652 18924
rect 22704 18952 22710 18964
rect 23198 18952 23204 18964
rect 22704 18924 23204 18952
rect 22704 18912 22710 18924
rect 23198 18912 23204 18924
rect 23256 18912 23262 18964
rect 26786 18912 26792 18964
rect 26844 18952 26850 18964
rect 32858 18952 32864 18964
rect 26844 18924 32864 18952
rect 26844 18912 26850 18924
rect 32858 18912 32864 18924
rect 32916 18912 32922 18964
rect 32953 18955 33011 18961
rect 32953 18921 32965 18955
rect 32999 18952 33011 18955
rect 34422 18952 34428 18964
rect 32999 18924 34428 18952
rect 32999 18921 33011 18924
rect 32953 18915 33011 18921
rect 34422 18912 34428 18924
rect 34480 18912 34486 18964
rect 19996 18884 20024 18912
rect 19306 18856 20024 18884
rect 20180 18884 20208 18912
rect 22005 18887 22063 18893
rect 20180 18856 21588 18884
rect 18616 18816 18644 18844
rect 14568 18788 18644 18816
rect 14568 18757 14596 18788
rect 19334 18776 19340 18828
rect 19392 18776 19398 18828
rect 19536 18788 19774 18816
rect 19536 18760 19564 18788
rect 14369 18751 14427 18757
rect 14369 18717 14381 18751
rect 14415 18717 14427 18751
rect 14369 18711 14427 18717
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18717 14611 18751
rect 14553 18711 14611 18717
rect 16758 18708 16764 18760
rect 16816 18708 16822 18760
rect 17678 18708 17684 18760
rect 17736 18708 17742 18760
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 12526 18640 12532 18692
rect 12584 18680 12590 18692
rect 13354 18680 13360 18692
rect 12584 18652 13360 18680
rect 12584 18640 12590 18652
rect 13354 18640 13360 18652
rect 13412 18680 13418 18692
rect 16776 18680 16804 18708
rect 17126 18680 17132 18692
rect 13412 18652 15516 18680
rect 16776 18652 17132 18680
rect 13412 18640 13418 18652
rect 15488 18624 15516 18652
rect 17126 18640 17132 18652
rect 17184 18680 17190 18692
rect 17972 18680 18000 18711
rect 18046 18708 18052 18760
rect 18104 18708 18110 18760
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18748 18291 18751
rect 18279 18720 18368 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 18340 18689 18368 18720
rect 18414 18708 18420 18760
rect 18472 18748 18478 18760
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 18472 18720 18521 18748
rect 18472 18708 18478 18720
rect 18509 18717 18521 18720
rect 18555 18717 18567 18751
rect 18509 18711 18567 18717
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18748 18659 18751
rect 18647 18720 18828 18748
rect 18647 18717 18659 18720
rect 18601 18711 18659 18717
rect 17184 18652 18000 18680
rect 18325 18683 18383 18689
rect 17184 18640 17190 18652
rect 18325 18649 18337 18683
rect 18371 18680 18383 18683
rect 18690 18680 18696 18692
rect 18371 18652 18696 18680
rect 18371 18649 18383 18652
rect 18325 18643 18383 18649
rect 18690 18640 18696 18652
rect 18748 18640 18754 18692
rect 18800 18680 18828 18720
rect 19242 18708 19248 18760
rect 19300 18708 19306 18760
rect 19518 18708 19524 18760
rect 19576 18708 19582 18760
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 19629 18680 19657 18708
rect 18800 18652 19657 18680
rect 19746 18680 19774 18788
rect 19978 18776 19984 18828
rect 20036 18776 20042 18828
rect 20165 18819 20223 18825
rect 20165 18785 20177 18819
rect 20211 18785 20223 18819
rect 20165 18779 20223 18785
rect 20441 18819 20499 18825
rect 20441 18785 20453 18819
rect 20487 18816 20499 18819
rect 20487 18788 20668 18816
rect 20487 18785 20499 18788
rect 20441 18779 20499 18785
rect 20180 18680 20208 18779
rect 20640 18760 20668 18788
rect 20533 18751 20591 18757
rect 20533 18717 20545 18751
rect 20579 18717 20591 18751
rect 20533 18711 20591 18717
rect 19746 18652 20208 18680
rect 18800 18624 18828 18652
rect 11388 18584 12204 18612
rect 11388 18572 11394 18584
rect 14182 18572 14188 18624
rect 14240 18572 14246 18624
rect 15470 18572 15476 18624
rect 15528 18572 15534 18624
rect 15746 18572 15752 18624
rect 15804 18612 15810 18624
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 15804 18584 17509 18612
rect 15804 18572 15810 18584
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 17497 18575 17555 18581
rect 18046 18572 18052 18624
rect 18104 18572 18110 18624
rect 18782 18572 18788 18624
rect 18840 18572 18846 18624
rect 18874 18572 18880 18624
rect 18932 18612 18938 18624
rect 20548 18612 20576 18711
rect 20622 18708 20628 18760
rect 20680 18708 20686 18760
rect 21560 18757 21588 18856
rect 22005 18853 22017 18887
rect 22051 18884 22063 18887
rect 25866 18884 25872 18896
rect 22051 18856 25872 18884
rect 22051 18853 22063 18856
rect 22005 18847 22063 18853
rect 25866 18844 25872 18856
rect 25924 18844 25930 18896
rect 27430 18844 27436 18896
rect 27488 18884 27494 18896
rect 33597 18887 33655 18893
rect 33597 18884 33609 18887
rect 27488 18856 33609 18884
rect 27488 18844 27494 18856
rect 33597 18853 33609 18856
rect 33643 18853 33655 18887
rect 33597 18847 33655 18853
rect 21821 18819 21879 18825
rect 21821 18785 21833 18819
rect 21867 18816 21879 18819
rect 22649 18819 22707 18825
rect 22649 18816 22661 18819
rect 21867 18788 22661 18816
rect 21867 18785 21879 18788
rect 21821 18779 21879 18785
rect 22649 18785 22661 18788
rect 22695 18816 22707 18819
rect 23474 18816 23480 18828
rect 22695 18788 23480 18816
rect 22695 18785 22707 18788
rect 22649 18779 22707 18785
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 33134 18816 33140 18828
rect 31036 18788 31616 18816
rect 21545 18751 21603 18757
rect 21545 18717 21557 18751
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 21634 18708 21640 18760
rect 21692 18708 21698 18760
rect 22370 18708 22376 18760
rect 22428 18708 22434 18760
rect 31036 18757 31064 18788
rect 31021 18751 31079 18757
rect 31021 18717 31033 18751
rect 31067 18717 31079 18751
rect 31021 18711 31079 18717
rect 31205 18751 31263 18757
rect 31205 18717 31217 18751
rect 31251 18748 31263 18751
rect 31294 18748 31300 18760
rect 31251 18720 31300 18748
rect 31251 18717 31263 18720
rect 31205 18711 31263 18717
rect 21174 18640 21180 18692
rect 21232 18640 21238 18692
rect 31036 18624 31064 18711
rect 31294 18708 31300 18720
rect 31352 18708 31358 18760
rect 31386 18708 31392 18760
rect 31444 18708 31450 18760
rect 31588 18757 31616 18788
rect 32508 18788 33140 18816
rect 32508 18757 32536 18788
rect 33134 18776 33140 18788
rect 33192 18776 33198 18828
rect 35434 18816 35440 18828
rect 34716 18788 35440 18816
rect 31573 18751 31631 18757
rect 31573 18717 31585 18751
rect 31619 18717 31631 18751
rect 31573 18711 31631 18717
rect 32401 18751 32459 18757
rect 32401 18717 32413 18751
rect 32447 18717 32459 18751
rect 32401 18711 32459 18717
rect 32493 18751 32551 18757
rect 32493 18717 32505 18751
rect 32539 18717 32551 18751
rect 32493 18711 32551 18717
rect 31481 18683 31539 18689
rect 31481 18649 31493 18683
rect 31527 18680 31539 18683
rect 32416 18680 32444 18711
rect 32674 18708 32680 18760
rect 32732 18708 32738 18760
rect 32766 18708 32772 18760
rect 32824 18708 32830 18760
rect 32950 18708 32956 18760
rect 33008 18748 33014 18760
rect 33689 18751 33747 18757
rect 33008 18720 33272 18748
rect 33008 18708 33014 18720
rect 33244 18680 33272 18720
rect 33689 18717 33701 18751
rect 33735 18748 33747 18751
rect 33962 18748 33968 18760
rect 33735 18720 33968 18748
rect 33735 18717 33747 18720
rect 33689 18711 33747 18717
rect 33962 18708 33968 18720
rect 34020 18708 34026 18760
rect 34716 18689 34744 18788
rect 35434 18776 35440 18788
rect 35492 18776 35498 18828
rect 36722 18776 36728 18828
rect 36780 18776 36786 18828
rect 34977 18751 35035 18757
rect 34977 18717 34989 18751
rect 35023 18748 35035 18751
rect 36909 18751 36967 18757
rect 36909 18748 36921 18751
rect 35023 18720 35204 18748
rect 35023 18717 35035 18720
rect 34977 18711 35035 18717
rect 34701 18683 34759 18689
rect 34701 18680 34713 18683
rect 31527 18652 33180 18680
rect 33244 18652 34713 18680
rect 31527 18649 31539 18652
rect 31481 18643 31539 18649
rect 33152 18624 33180 18652
rect 34701 18649 34713 18652
rect 34747 18649 34759 18683
rect 34701 18643 34759 18649
rect 35176 18624 35204 18720
rect 36832 18720 36921 18748
rect 36832 18692 36860 18720
rect 36909 18717 36921 18720
rect 36955 18717 36967 18751
rect 36909 18711 36967 18717
rect 36814 18640 36820 18692
rect 36872 18640 36878 18692
rect 20990 18621 20996 18624
rect 18932 18584 20576 18612
rect 20977 18615 20996 18621
rect 18932 18572 18938 18584
rect 20977 18581 20989 18615
rect 20977 18575 20996 18581
rect 20990 18572 20996 18575
rect 21048 18572 21054 18624
rect 22186 18572 22192 18624
rect 22244 18572 22250 18624
rect 25590 18572 25596 18624
rect 25648 18612 25654 18624
rect 26050 18612 26056 18624
rect 25648 18584 26056 18612
rect 25648 18572 25654 18584
rect 26050 18572 26056 18584
rect 26108 18612 26114 18624
rect 28442 18612 28448 18624
rect 26108 18584 28448 18612
rect 26108 18572 26114 18584
rect 28442 18572 28448 18584
rect 28500 18612 28506 18624
rect 30742 18612 30748 18624
rect 28500 18584 30748 18612
rect 28500 18572 28506 18584
rect 30742 18572 30748 18584
rect 30800 18572 30806 18624
rect 31018 18572 31024 18624
rect 31076 18572 31082 18624
rect 31202 18572 31208 18624
rect 31260 18572 31266 18624
rect 32306 18572 32312 18624
rect 32364 18612 32370 18624
rect 32950 18612 32956 18624
rect 32364 18584 32956 18612
rect 32364 18572 32370 18584
rect 32950 18572 32956 18584
rect 33008 18572 33014 18624
rect 33134 18572 33140 18624
rect 33192 18572 33198 18624
rect 34790 18572 34796 18624
rect 34848 18621 34854 18624
rect 34848 18575 34857 18621
rect 34885 18615 34943 18621
rect 34885 18581 34897 18615
rect 34931 18612 34943 18615
rect 34974 18612 34980 18624
rect 34931 18584 34980 18612
rect 34931 18581 34943 18584
rect 34885 18575 34943 18581
rect 34848 18572 34854 18575
rect 34974 18572 34980 18584
rect 35032 18572 35038 18624
rect 35158 18572 35164 18624
rect 35216 18572 35222 18624
rect 37090 18572 37096 18624
rect 37148 18572 37154 18624
rect 1104 18522 38272 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38272 18522
rect 1104 18448 38272 18470
rect 4246 18408 4252 18420
rect 2332 18380 4252 18408
rect 2332 18281 2360 18380
rect 4246 18368 4252 18380
rect 4304 18368 4310 18420
rect 13814 18408 13820 18420
rect 4356 18380 9536 18408
rect 4356 18349 4384 18380
rect 4341 18343 4399 18349
rect 4341 18309 4353 18343
rect 4387 18309 4399 18343
rect 4341 18303 4399 18309
rect 8294 18300 8300 18352
rect 8352 18300 8358 18352
rect 9508 18349 9536 18380
rect 11256 18380 13820 18408
rect 9493 18343 9551 18349
rect 9493 18309 9505 18343
rect 9539 18340 9551 18343
rect 10226 18340 10232 18352
rect 9539 18312 10232 18340
rect 9539 18309 9551 18312
rect 9493 18303 9551 18309
rect 10226 18300 10232 18312
rect 10284 18300 10290 18352
rect 10778 18300 10784 18352
rect 10836 18340 10842 18352
rect 11256 18349 11284 18380
rect 13814 18368 13820 18380
rect 13872 18368 13878 18420
rect 13906 18368 13912 18420
rect 13964 18368 13970 18420
rect 14182 18368 14188 18420
rect 14240 18368 14246 18420
rect 15378 18368 15384 18420
rect 15436 18368 15442 18420
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 19429 18411 19487 18417
rect 19429 18408 19441 18411
rect 19392 18380 19441 18408
rect 19392 18368 19398 18380
rect 19429 18377 19441 18380
rect 19475 18377 19487 18411
rect 22094 18408 22100 18420
rect 19429 18371 19487 18377
rect 19536 18380 22100 18408
rect 11241 18343 11299 18349
rect 11241 18340 11253 18343
rect 10836 18312 11253 18340
rect 10836 18300 10842 18312
rect 11241 18309 11253 18312
rect 11287 18309 11299 18343
rect 11241 18303 11299 18309
rect 11330 18300 11336 18352
rect 11388 18300 11394 18352
rect 12069 18343 12127 18349
rect 12069 18309 12081 18343
rect 12115 18340 12127 18343
rect 12250 18340 12256 18352
rect 12115 18312 12256 18340
rect 12115 18309 12127 18312
rect 12069 18303 12127 18309
rect 12250 18300 12256 18312
rect 12308 18300 12314 18352
rect 14200 18340 14228 18368
rect 14200 18312 14504 18340
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18272 1915 18275
rect 2317 18275 2375 18281
rect 1903 18244 2268 18272
rect 1903 18241 1915 18244
rect 1857 18235 1915 18241
rect 1670 18164 1676 18216
rect 1728 18204 1734 18216
rect 2133 18207 2191 18213
rect 2133 18204 2145 18207
rect 1728 18176 2145 18204
rect 1728 18164 1734 18176
rect 2133 18173 2145 18176
rect 2179 18173 2191 18207
rect 2240 18204 2268 18244
rect 2317 18241 2329 18275
rect 2363 18241 2375 18275
rect 2317 18235 2375 18241
rect 6181 18275 6239 18281
rect 6181 18241 6193 18275
rect 6227 18272 6239 18275
rect 6730 18272 6736 18284
rect 6227 18244 6736 18272
rect 6227 18241 6239 18244
rect 6181 18235 6239 18241
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 11348 18272 11376 18300
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 11348 18244 11529 18272
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 11517 18235 11575 18241
rect 11698 18232 11704 18284
rect 11756 18232 11762 18284
rect 12342 18232 12348 18284
rect 12400 18232 12406 18284
rect 12526 18232 12532 18284
rect 12584 18232 12590 18284
rect 12802 18232 12808 18284
rect 12860 18272 12866 18284
rect 13998 18272 14004 18284
rect 12860 18244 14004 18272
rect 12860 18232 12866 18244
rect 13998 18232 14004 18244
rect 14056 18272 14062 18284
rect 14093 18275 14151 18281
rect 14093 18272 14105 18275
rect 14056 18244 14105 18272
rect 14056 18232 14062 18244
rect 14093 18241 14105 18244
rect 14139 18241 14151 18275
rect 14093 18235 14151 18241
rect 14182 18232 14188 18284
rect 14240 18272 14246 18284
rect 14476 18281 14504 18312
rect 16850 18300 16856 18352
rect 16908 18340 16914 18352
rect 17586 18340 17592 18352
rect 16908 18312 17592 18340
rect 16908 18300 16914 18312
rect 14277 18275 14335 18281
rect 14277 18272 14289 18275
rect 14240 18244 14289 18272
rect 14240 18232 14246 18244
rect 14277 18241 14289 18244
rect 14323 18241 14335 18275
rect 14277 18235 14335 18241
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 16390 18232 16396 18284
rect 16448 18272 16454 18284
rect 16945 18275 17003 18281
rect 16945 18272 16957 18275
rect 16448 18244 16957 18272
rect 16448 18232 16454 18244
rect 16945 18241 16957 18244
rect 16991 18272 17003 18275
rect 17034 18272 17040 18284
rect 16991 18244 17040 18272
rect 16991 18241 17003 18244
rect 16945 18235 17003 18241
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 17144 18281 17172 18312
rect 17586 18300 17592 18312
rect 17644 18300 17650 18352
rect 18414 18300 18420 18352
rect 18472 18340 18478 18352
rect 18472 18312 18920 18340
rect 18472 18300 18478 18312
rect 17129 18275 17187 18281
rect 17129 18241 17141 18275
rect 17175 18241 17187 18275
rect 17129 18235 17187 18241
rect 18230 18232 18236 18284
rect 18288 18272 18294 18284
rect 18892 18281 18920 18312
rect 19058 18300 19064 18352
rect 19116 18340 19122 18352
rect 19536 18340 19564 18380
rect 22094 18368 22100 18380
rect 22152 18368 22158 18420
rect 25593 18411 25651 18417
rect 25593 18377 25605 18411
rect 25639 18408 25651 18411
rect 25639 18380 30696 18408
rect 25639 18377 25651 18380
rect 25593 18371 25651 18377
rect 19116 18312 19564 18340
rect 19889 18343 19947 18349
rect 19116 18300 19122 18312
rect 19889 18309 19901 18343
rect 19935 18340 19947 18343
rect 19978 18340 19984 18352
rect 19935 18312 19984 18340
rect 19935 18309 19947 18312
rect 19889 18303 19947 18309
rect 19978 18300 19984 18312
rect 20036 18300 20042 18352
rect 22646 18340 22652 18352
rect 22480 18312 22652 18340
rect 18785 18275 18843 18281
rect 18785 18272 18797 18275
rect 18288 18244 18797 18272
rect 18288 18232 18294 18244
rect 18785 18241 18797 18244
rect 18831 18241 18843 18275
rect 18785 18235 18843 18241
rect 18877 18275 18935 18281
rect 18877 18241 18889 18275
rect 18923 18241 18935 18275
rect 18877 18235 18935 18241
rect 4062 18204 4068 18216
rect 2240 18176 4068 18204
rect 2133 18167 2191 18173
rect 2148 18136 2176 18167
rect 4062 18164 4068 18176
rect 4120 18164 4126 18216
rect 5902 18164 5908 18216
rect 5960 18164 5966 18216
rect 6638 18204 6644 18216
rect 6196 18176 6644 18204
rect 3694 18136 3700 18148
rect 2148 18108 3700 18136
rect 3694 18096 3700 18108
rect 3752 18096 3758 18148
rect 6196 18080 6224 18176
rect 6638 18164 6644 18176
rect 6696 18204 6702 18216
rect 7561 18207 7619 18213
rect 7561 18204 7573 18207
rect 6696 18176 7573 18204
rect 6696 18164 6702 18176
rect 7561 18173 7573 18176
rect 7607 18173 7619 18207
rect 7561 18167 7619 18173
rect 7837 18207 7895 18213
rect 7837 18173 7849 18207
rect 7883 18204 7895 18207
rect 7926 18204 7932 18216
rect 7883 18176 7932 18204
rect 7883 18173 7895 18176
rect 7837 18167 7895 18173
rect 2038 18028 2044 18080
rect 2096 18028 2102 18080
rect 2498 18028 2504 18080
rect 2556 18028 2562 18080
rect 2958 18028 2964 18080
rect 3016 18068 3022 18080
rect 3053 18071 3111 18077
rect 3053 18068 3065 18071
rect 3016 18040 3065 18068
rect 3016 18028 3022 18040
rect 3053 18037 3065 18040
rect 3099 18068 3111 18071
rect 3510 18068 3516 18080
rect 3099 18040 3516 18068
rect 3099 18037 3111 18040
rect 3053 18031 3111 18037
rect 3510 18028 3516 18040
rect 3568 18028 3574 18080
rect 6178 18028 6184 18080
rect 6236 18028 6242 18080
rect 7576 18068 7604 18167
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 9214 18164 9220 18216
rect 9272 18204 9278 18216
rect 9272 18176 12020 18204
rect 9272 18164 9278 18176
rect 10778 18136 10784 18148
rect 8864 18108 10784 18136
rect 8864 18080 8892 18108
rect 10778 18096 10784 18108
rect 10836 18096 10842 18148
rect 11146 18096 11152 18148
rect 11204 18136 11210 18148
rect 11701 18139 11759 18145
rect 11701 18136 11713 18139
rect 11204 18108 11713 18136
rect 11204 18096 11210 18108
rect 11701 18105 11713 18108
rect 11747 18105 11759 18139
rect 11992 18136 12020 18176
rect 12066 18164 12072 18216
rect 12124 18204 12130 18216
rect 12161 18207 12219 18213
rect 12161 18204 12173 18207
rect 12124 18176 12173 18204
rect 12124 18164 12130 18176
rect 12161 18173 12173 18176
rect 12207 18173 12219 18207
rect 12161 18167 12219 18173
rect 12710 18164 12716 18216
rect 12768 18204 12774 18216
rect 13906 18204 13912 18216
rect 12768 18176 13912 18204
rect 12768 18164 12774 18176
rect 13906 18164 13912 18176
rect 13964 18204 13970 18216
rect 14734 18204 14740 18216
rect 13964 18176 14740 18204
rect 13964 18164 13970 18176
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 15562 18164 15568 18216
rect 15620 18164 15626 18216
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18173 15715 18207
rect 15657 18167 15715 18173
rect 12728 18136 12756 18164
rect 11992 18108 12756 18136
rect 11701 18099 11759 18105
rect 15470 18096 15476 18148
rect 15528 18136 15534 18148
rect 15672 18136 15700 18167
rect 15930 18164 15936 18216
rect 15988 18204 15994 18216
rect 16025 18207 16083 18213
rect 16025 18204 16037 18207
rect 15988 18176 16037 18204
rect 15988 18164 15994 18176
rect 16025 18173 16037 18176
rect 16071 18173 16083 18207
rect 18892 18204 18920 18235
rect 18966 18232 18972 18284
rect 19024 18272 19030 18284
rect 19245 18275 19303 18281
rect 19245 18272 19257 18275
rect 19024 18244 19257 18272
rect 19024 18232 19030 18244
rect 19245 18241 19257 18244
rect 19291 18241 19303 18275
rect 19245 18235 19303 18241
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 19426 18204 19432 18216
rect 18892 18176 19432 18204
rect 16025 18167 16083 18173
rect 19426 18164 19432 18176
rect 19484 18164 19490 18216
rect 19536 18136 19564 18235
rect 19610 18232 19616 18284
rect 19668 18232 19674 18284
rect 20438 18232 20444 18284
rect 20496 18232 20502 18284
rect 22370 18232 22376 18284
rect 22428 18232 22434 18284
rect 22480 18281 22508 18312
rect 22646 18300 22652 18312
rect 22704 18300 22710 18352
rect 29454 18300 29460 18352
rect 29512 18340 29518 18352
rect 30374 18340 30380 18352
rect 29512 18312 30380 18340
rect 29512 18300 29518 18312
rect 22465 18275 22523 18281
rect 22465 18241 22477 18275
rect 22511 18241 22523 18275
rect 22465 18235 22523 18241
rect 22554 18232 22560 18284
rect 22612 18272 22618 18284
rect 22741 18275 22799 18281
rect 22741 18272 22753 18275
rect 22612 18244 22753 18272
rect 22612 18232 22618 18244
rect 22741 18241 22753 18244
rect 22787 18241 22799 18275
rect 22741 18235 22799 18241
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18272 23351 18275
rect 23934 18272 23940 18284
rect 23339 18244 23940 18272
rect 23339 18241 23351 18244
rect 23293 18235 23351 18241
rect 23934 18232 23940 18244
rect 23992 18232 23998 18284
rect 25038 18232 25044 18284
rect 25096 18232 25102 18284
rect 25130 18232 25136 18284
rect 25188 18272 25194 18284
rect 25225 18275 25283 18281
rect 25225 18272 25237 18275
rect 25188 18244 25237 18272
rect 25188 18232 25194 18244
rect 25225 18241 25237 18244
rect 25271 18241 25283 18275
rect 25225 18235 25283 18241
rect 25317 18275 25375 18281
rect 25317 18241 25329 18275
rect 25363 18241 25375 18275
rect 25317 18235 25375 18241
rect 20456 18136 20484 18232
rect 22388 18204 22416 18232
rect 22925 18207 22983 18213
rect 22925 18204 22937 18207
rect 22388 18176 22937 18204
rect 22925 18173 22937 18176
rect 22971 18173 22983 18207
rect 22925 18167 22983 18173
rect 23658 18164 23664 18216
rect 23716 18204 23722 18216
rect 25332 18204 25360 18235
rect 25406 18232 25412 18284
rect 25464 18232 25470 18284
rect 25869 18275 25927 18281
rect 25869 18241 25881 18275
rect 25915 18272 25927 18275
rect 26050 18272 26056 18284
rect 25915 18244 26056 18272
rect 25915 18241 25927 18244
rect 25869 18235 25927 18241
rect 26050 18232 26056 18244
rect 26108 18232 26114 18284
rect 27982 18232 27988 18284
rect 28040 18232 28046 18284
rect 28166 18232 28172 18284
rect 28224 18232 28230 18284
rect 29564 18281 29592 18312
rect 30116 18281 30144 18312
rect 30374 18300 30380 18312
rect 30432 18300 30438 18352
rect 30668 18340 30696 18380
rect 31202 18368 31208 18420
rect 31260 18408 31266 18420
rect 31260 18380 31754 18408
rect 31260 18368 31266 18380
rect 30668 18312 30972 18340
rect 29549 18275 29607 18281
rect 29549 18241 29561 18275
rect 29595 18241 29607 18275
rect 29549 18235 29607 18241
rect 29733 18275 29791 18281
rect 29733 18241 29745 18275
rect 29779 18272 29791 18275
rect 30101 18275 30159 18281
rect 29779 18244 29868 18272
rect 29779 18241 29791 18244
rect 29733 18235 29791 18241
rect 23716 18176 25360 18204
rect 23716 18164 23722 18176
rect 25774 18164 25780 18216
rect 25832 18164 25838 18216
rect 28184 18204 28212 18232
rect 28626 18204 28632 18216
rect 28184 18176 28632 18204
rect 28626 18164 28632 18176
rect 28684 18164 28690 18216
rect 15528 18108 20484 18136
rect 23569 18139 23627 18145
rect 15528 18096 15534 18108
rect 23569 18105 23581 18139
rect 23615 18105 23627 18139
rect 23569 18099 23627 18105
rect 8846 18068 8852 18080
rect 7576 18040 8852 18068
rect 8846 18028 8852 18040
rect 8904 18028 8910 18080
rect 9122 18028 9128 18080
rect 9180 18068 9186 18080
rect 9309 18071 9367 18077
rect 9309 18068 9321 18071
rect 9180 18040 9321 18068
rect 9180 18028 9186 18040
rect 9309 18037 9321 18040
rect 9355 18037 9367 18071
rect 9309 18031 9367 18037
rect 14274 18028 14280 18080
rect 14332 18068 14338 18080
rect 14642 18068 14648 18080
rect 14332 18040 14648 18068
rect 14332 18028 14338 18040
rect 14642 18028 14648 18040
rect 14700 18028 14706 18080
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 16942 18068 16948 18080
rect 15436 18040 16948 18068
rect 15436 18028 15442 18040
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 17954 18028 17960 18080
rect 18012 18068 18018 18080
rect 18417 18071 18475 18077
rect 18417 18068 18429 18071
rect 18012 18040 18429 18068
rect 18012 18028 18018 18040
rect 18417 18037 18429 18040
rect 18463 18068 18475 18071
rect 18506 18068 18512 18080
rect 18463 18040 18512 18068
rect 18463 18037 18475 18040
rect 18417 18031 18475 18037
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 18874 18028 18880 18080
rect 18932 18068 18938 18080
rect 19153 18071 19211 18077
rect 19153 18068 19165 18071
rect 18932 18040 19165 18068
rect 18932 18028 18938 18040
rect 19153 18037 19165 18040
rect 19199 18037 19211 18071
rect 19153 18031 19211 18037
rect 19242 18028 19248 18080
rect 19300 18068 19306 18080
rect 19610 18068 19616 18080
rect 19300 18040 19616 18068
rect 19300 18028 19306 18040
rect 19610 18028 19616 18040
rect 19668 18028 19674 18080
rect 23584 18068 23612 18099
rect 24670 18096 24676 18148
rect 24728 18136 24734 18148
rect 25682 18136 25688 18148
rect 24728 18108 25688 18136
rect 24728 18096 24734 18108
rect 25682 18096 25688 18108
rect 25740 18096 25746 18148
rect 26234 18096 26240 18148
rect 26292 18096 26298 18148
rect 28902 18096 28908 18148
rect 28960 18136 28966 18148
rect 29840 18136 29868 18244
rect 30101 18241 30113 18275
rect 30147 18241 30159 18275
rect 30653 18275 30711 18281
rect 30653 18272 30665 18275
rect 30101 18235 30159 18241
rect 30208 18244 30665 18272
rect 29914 18164 29920 18216
rect 29972 18204 29978 18216
rect 30208 18204 30236 18244
rect 30653 18241 30665 18244
rect 30699 18272 30711 18275
rect 30834 18272 30840 18284
rect 30699 18244 30840 18272
rect 30699 18241 30711 18244
rect 30653 18235 30711 18241
rect 30834 18232 30840 18244
rect 30892 18232 30898 18284
rect 30944 18272 30972 18312
rect 31294 18300 31300 18352
rect 31352 18300 31358 18352
rect 31726 18340 31754 18380
rect 32674 18368 32680 18420
rect 32732 18368 32738 18420
rect 32769 18411 32827 18417
rect 32769 18377 32781 18411
rect 32815 18408 32827 18411
rect 34146 18408 34152 18420
rect 32815 18380 34152 18408
rect 32815 18377 32827 18380
rect 32769 18371 32827 18377
rect 34146 18368 34152 18380
rect 34204 18408 34210 18420
rect 34241 18411 34299 18417
rect 34241 18408 34253 18411
rect 34204 18380 34253 18408
rect 34204 18368 34210 18380
rect 34241 18377 34253 18380
rect 34287 18377 34299 18411
rect 34241 18371 34299 18377
rect 34790 18368 34796 18420
rect 34848 18368 34854 18420
rect 37090 18368 37096 18420
rect 37148 18368 37154 18420
rect 32125 18343 32183 18349
rect 32125 18340 32137 18343
rect 31680 18312 32137 18340
rect 31018 18272 31024 18284
rect 30944 18244 31024 18272
rect 31018 18232 31024 18244
rect 31076 18232 31082 18284
rect 31205 18275 31263 18281
rect 31205 18241 31217 18275
rect 31251 18272 31263 18275
rect 31312 18272 31340 18300
rect 31680 18281 31708 18312
rect 32125 18309 32137 18312
rect 32171 18309 32183 18343
rect 32692 18340 32720 18368
rect 32953 18343 33011 18349
rect 32953 18340 32965 18343
rect 32125 18303 32183 18309
rect 32232 18312 32965 18340
rect 31251 18244 31340 18272
rect 31389 18275 31447 18281
rect 31251 18241 31263 18244
rect 31205 18235 31263 18241
rect 31389 18241 31401 18275
rect 31435 18272 31447 18275
rect 31481 18275 31539 18281
rect 31481 18272 31493 18275
rect 31435 18244 31493 18272
rect 31435 18241 31447 18244
rect 31389 18235 31447 18241
rect 31481 18241 31493 18244
rect 31527 18241 31539 18275
rect 31481 18235 31539 18241
rect 31665 18275 31723 18281
rect 31665 18241 31677 18275
rect 31711 18241 31723 18275
rect 31665 18235 31723 18241
rect 31849 18275 31907 18281
rect 31849 18241 31861 18275
rect 31895 18272 31907 18275
rect 32030 18272 32036 18284
rect 31895 18244 32036 18272
rect 31895 18241 31907 18244
rect 31849 18235 31907 18241
rect 32030 18232 32036 18244
rect 32088 18272 32094 18284
rect 32232 18272 32260 18312
rect 32953 18309 32965 18312
rect 32999 18309 33011 18343
rect 32953 18303 33011 18309
rect 33134 18300 33140 18352
rect 33192 18300 33198 18352
rect 34072 18312 34744 18340
rect 32088 18244 32260 18272
rect 32088 18232 32094 18244
rect 32674 18232 32680 18284
rect 32732 18272 32738 18284
rect 32861 18275 32919 18281
rect 32861 18272 32873 18275
rect 32732 18244 32873 18272
rect 32732 18232 32738 18244
rect 32861 18241 32873 18244
rect 32907 18241 32919 18275
rect 32861 18235 32919 18241
rect 29972 18176 30236 18204
rect 30469 18207 30527 18213
rect 29972 18164 29978 18176
rect 30469 18173 30481 18207
rect 30515 18204 30527 18207
rect 31570 18204 31576 18216
rect 30515 18176 31576 18204
rect 30515 18173 30527 18176
rect 30469 18167 30527 18173
rect 31570 18164 31576 18176
rect 31628 18164 31634 18216
rect 32490 18164 32496 18216
rect 32548 18164 32554 18216
rect 32582 18164 32588 18216
rect 32640 18164 32646 18216
rect 34072 18213 34100 18312
rect 34333 18275 34391 18281
rect 34333 18241 34345 18275
rect 34379 18241 34391 18275
rect 34333 18235 34391 18241
rect 34057 18207 34115 18213
rect 34057 18204 34069 18207
rect 33060 18176 34069 18204
rect 32122 18136 32128 18148
rect 28960 18108 32128 18136
rect 28960 18096 28966 18108
rect 32122 18096 32128 18108
rect 32180 18136 32186 18148
rect 32766 18136 32772 18148
rect 32180 18108 32772 18136
rect 32180 18096 32186 18108
rect 32766 18096 32772 18108
rect 32824 18096 32830 18148
rect 26510 18068 26516 18080
rect 23584 18040 26516 18068
rect 26510 18028 26516 18040
rect 26568 18028 26574 18080
rect 27890 18028 27896 18080
rect 27948 18068 27954 18080
rect 28077 18071 28135 18077
rect 28077 18068 28089 18071
rect 27948 18040 28089 18068
rect 27948 18028 27954 18040
rect 28077 18037 28089 18040
rect 28123 18037 28135 18071
rect 28077 18031 28135 18037
rect 29546 18028 29552 18080
rect 29604 18068 29610 18080
rect 29914 18068 29920 18080
rect 29604 18040 29920 18068
rect 29604 18028 29610 18040
rect 29914 18028 29920 18040
rect 29972 18028 29978 18080
rect 31754 18028 31760 18080
rect 31812 18068 31818 18080
rect 33060 18068 33088 18176
rect 34057 18173 34069 18176
rect 34103 18173 34115 18207
rect 34057 18167 34115 18173
rect 33137 18139 33195 18145
rect 33137 18105 33149 18139
rect 33183 18136 33195 18139
rect 34348 18136 34376 18235
rect 34716 18204 34744 18312
rect 34808 18281 34836 18368
rect 35618 18340 35624 18352
rect 35084 18312 35624 18340
rect 34793 18275 34851 18281
rect 34793 18241 34805 18275
rect 34839 18241 34851 18275
rect 34793 18235 34851 18241
rect 34974 18232 34980 18284
rect 35032 18232 35038 18284
rect 35084 18204 35112 18312
rect 35618 18300 35624 18312
rect 35676 18300 35682 18352
rect 35158 18232 35164 18284
rect 35216 18232 35222 18284
rect 36909 18275 36967 18281
rect 36909 18241 36921 18275
rect 36955 18272 36967 18275
rect 37108 18272 37136 18368
rect 37182 18300 37188 18352
rect 37240 18340 37246 18352
rect 37240 18312 37596 18340
rect 37240 18300 37246 18312
rect 37568 18281 37596 18312
rect 36955 18244 37136 18272
rect 37553 18275 37611 18281
rect 36955 18241 36967 18244
rect 36909 18235 36967 18241
rect 37553 18241 37565 18275
rect 37599 18241 37611 18275
rect 37553 18235 37611 18241
rect 34716 18176 35112 18204
rect 33183 18108 34376 18136
rect 34701 18139 34759 18145
rect 33183 18105 33195 18108
rect 33137 18099 33195 18105
rect 34701 18105 34713 18139
rect 34747 18136 34759 18139
rect 35176 18136 35204 18232
rect 34747 18108 35204 18136
rect 34747 18105 34759 18108
rect 34701 18099 34759 18105
rect 31812 18040 33088 18068
rect 31812 18028 31818 18040
rect 33962 18028 33968 18080
rect 34020 18068 34026 18080
rect 34885 18071 34943 18077
rect 34885 18068 34897 18071
rect 34020 18040 34897 18068
rect 34020 18028 34026 18040
rect 34885 18037 34897 18040
rect 34931 18037 34943 18071
rect 34885 18031 34943 18037
rect 37093 18071 37151 18077
rect 37093 18037 37105 18071
rect 37139 18068 37151 18071
rect 37550 18068 37556 18080
rect 37139 18040 37556 18068
rect 37139 18037 37151 18040
rect 37093 18031 37151 18037
rect 37550 18028 37556 18040
rect 37608 18028 37614 18080
rect 37829 18071 37887 18077
rect 37829 18037 37841 18071
rect 37875 18068 37887 18071
rect 37875 18040 38424 18068
rect 37875 18037 37887 18040
rect 37829 18031 37887 18037
rect 38396 18012 38424 18040
rect 1104 17978 38272 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38272 17978
rect 38378 17960 38384 18012
rect 38436 17960 38442 18012
rect 1104 17904 38272 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 2041 17867 2099 17873
rect 2041 17864 2053 17867
rect 1820 17836 2053 17864
rect 1820 17824 1826 17836
rect 2041 17833 2053 17836
rect 2087 17833 2099 17867
rect 2041 17827 2099 17833
rect 2130 17824 2136 17876
rect 2188 17864 2194 17876
rect 2961 17867 3019 17873
rect 2961 17864 2973 17867
rect 2188 17836 2973 17864
rect 2188 17824 2194 17836
rect 2961 17833 2973 17836
rect 3007 17833 3019 17867
rect 5626 17864 5632 17876
rect 2961 17827 3019 17833
rect 3344 17836 5632 17864
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17728 1639 17731
rect 1670 17728 1676 17740
rect 1627 17700 1676 17728
rect 1627 17697 1639 17700
rect 1581 17691 1639 17697
rect 1670 17688 1676 17700
rect 1728 17688 1734 17740
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 1946 17660 1952 17672
rect 1811 17632 1952 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 2038 17620 2044 17672
rect 2096 17660 2102 17672
rect 3344 17669 3372 17836
rect 5626 17824 5632 17836
rect 5684 17824 5690 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 6972 17836 7696 17864
rect 6972 17824 6978 17836
rect 7668 17796 7696 17836
rect 7742 17824 7748 17876
rect 7800 17864 7806 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 7800 17836 7849 17864
rect 7800 17824 7806 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 7837 17827 7895 17833
rect 7926 17824 7932 17876
rect 7984 17864 7990 17876
rect 8021 17867 8079 17873
rect 8021 17864 8033 17867
rect 7984 17836 8033 17864
rect 7984 17824 7990 17836
rect 8021 17833 8033 17836
rect 8067 17833 8079 17867
rect 9858 17864 9864 17876
rect 8021 17827 8079 17833
rect 8864 17836 9864 17864
rect 8294 17796 8300 17808
rect 7668 17768 8300 17796
rect 8294 17756 8300 17768
rect 8352 17756 8358 17808
rect 3510 17688 3516 17740
rect 3568 17728 3574 17740
rect 3970 17728 3976 17740
rect 3568 17700 3976 17728
rect 3568 17688 3574 17700
rect 3970 17688 3976 17700
rect 4028 17688 4034 17740
rect 5442 17688 5448 17740
rect 5500 17688 5506 17740
rect 8864 17728 8892 17836
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 11333 17867 11391 17873
rect 11333 17833 11345 17867
rect 11379 17864 11391 17867
rect 11698 17864 11704 17876
rect 11379 17836 11704 17864
rect 11379 17833 11391 17836
rect 11333 17827 11391 17833
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 12434 17864 12440 17876
rect 11808 17836 12440 17864
rect 8941 17799 8999 17805
rect 8941 17765 8953 17799
rect 8987 17765 8999 17799
rect 8941 17759 8999 17765
rect 11241 17799 11299 17805
rect 11241 17765 11253 17799
rect 11287 17796 11299 17799
rect 11808 17796 11836 17836
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 12526 17824 12532 17876
rect 12584 17864 12590 17876
rect 12805 17867 12863 17873
rect 12805 17864 12817 17867
rect 12584 17836 12817 17864
rect 12584 17824 12590 17836
rect 12805 17833 12817 17836
rect 12851 17833 12863 17867
rect 12805 17827 12863 17833
rect 13078 17824 13084 17876
rect 13136 17864 13142 17876
rect 14734 17864 14740 17876
rect 13136 17836 14740 17864
rect 13136 17824 13142 17836
rect 14734 17824 14740 17836
rect 14792 17824 14798 17876
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 15289 17867 15347 17873
rect 15289 17864 15301 17867
rect 15252 17836 15301 17864
rect 15252 17824 15258 17836
rect 15289 17833 15301 17836
rect 15335 17833 15347 17867
rect 20625 17867 20683 17873
rect 20625 17864 20637 17867
rect 15289 17827 15347 17833
rect 16500 17836 20637 17864
rect 12544 17796 12572 17824
rect 16025 17799 16083 17805
rect 16025 17796 16037 17799
rect 11287 17768 11836 17796
rect 12452 17768 12572 17796
rect 12636 17768 16037 17796
rect 11287 17765 11299 17768
rect 11241 17759 11299 17765
rect 5644 17700 8892 17728
rect 2225 17663 2283 17669
rect 2225 17660 2237 17663
rect 2096 17632 2237 17660
rect 2096 17620 2102 17632
rect 2225 17629 2237 17632
rect 2271 17629 2283 17663
rect 2225 17623 2283 17629
rect 3237 17663 3295 17669
rect 3237 17629 3249 17663
rect 3283 17629 3295 17663
rect 3237 17623 3295 17629
rect 3329 17663 3387 17669
rect 3329 17629 3341 17663
rect 3375 17629 3387 17663
rect 3329 17623 3387 17629
rect 1946 17484 1952 17536
rect 2004 17484 2010 17536
rect 3252 17524 3280 17623
rect 3418 17620 3424 17672
rect 3476 17620 3482 17672
rect 3605 17663 3663 17669
rect 3605 17629 3617 17663
rect 3651 17660 3663 17663
rect 3694 17660 3700 17672
rect 3651 17632 3700 17660
rect 3651 17629 3663 17632
rect 3605 17623 3663 17629
rect 3694 17620 3700 17632
rect 3752 17620 3758 17672
rect 5460 17660 5488 17688
rect 5382 17632 5488 17660
rect 4246 17552 4252 17604
rect 4304 17552 4310 17604
rect 5644 17524 5672 17700
rect 6089 17663 6147 17669
rect 6089 17629 6101 17663
rect 6135 17629 6147 17663
rect 6089 17623 6147 17629
rect 8205 17663 8263 17669
rect 8205 17629 8217 17663
rect 8251 17660 8263 17663
rect 8956 17660 8984 17759
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 9401 17731 9459 17737
rect 9401 17728 9413 17731
rect 9180 17700 9413 17728
rect 9180 17688 9186 17700
rect 9401 17697 9413 17700
rect 9447 17697 9459 17731
rect 9401 17691 9459 17697
rect 9493 17731 9551 17737
rect 9493 17697 9505 17731
rect 9539 17697 9551 17731
rect 9493 17691 9551 17697
rect 9508 17660 9536 17691
rect 10042 17688 10048 17740
rect 10100 17728 10106 17740
rect 10873 17731 10931 17737
rect 10100 17700 10548 17728
rect 10100 17688 10106 17700
rect 10520 17672 10548 17700
rect 10873 17697 10885 17731
rect 10919 17728 10931 17731
rect 11146 17728 11152 17740
rect 10919 17700 11152 17728
rect 10919 17697 10931 17700
rect 10873 17691 10931 17697
rect 11146 17688 11152 17700
rect 11204 17688 11210 17740
rect 11606 17688 11612 17740
rect 11664 17728 11670 17740
rect 11793 17731 11851 17737
rect 11793 17728 11805 17731
rect 11664 17700 11805 17728
rect 11664 17688 11670 17700
rect 11793 17697 11805 17700
rect 11839 17697 11851 17731
rect 11793 17691 11851 17697
rect 11974 17688 11980 17740
rect 12032 17688 12038 17740
rect 8251 17632 8984 17660
rect 9232 17632 9536 17660
rect 10137 17663 10195 17669
rect 8251 17629 8263 17632
rect 8205 17623 8263 17629
rect 6104 17592 6132 17623
rect 6104 17564 6224 17592
rect 6196 17536 6224 17564
rect 6362 17552 6368 17604
rect 6420 17552 6426 17604
rect 6914 17552 6920 17604
rect 6972 17552 6978 17604
rect 3252 17496 5672 17524
rect 5718 17484 5724 17536
rect 5776 17484 5782 17536
rect 6178 17484 6184 17536
rect 6236 17484 6242 17536
rect 7190 17484 7196 17536
rect 7248 17524 7254 17536
rect 7374 17524 7380 17536
rect 7248 17496 7380 17524
rect 7248 17484 7254 17496
rect 7374 17484 7380 17496
rect 7432 17524 7438 17536
rect 9232 17524 9260 17632
rect 10137 17629 10149 17663
rect 10183 17629 10195 17663
rect 10137 17623 10195 17629
rect 10152 17592 10180 17623
rect 10318 17620 10324 17672
rect 10376 17660 10382 17672
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 10376 17632 10425 17660
rect 10376 17620 10382 17632
rect 10413 17629 10425 17632
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 10502 17620 10508 17672
rect 10560 17620 10566 17672
rect 10594 17620 10600 17672
rect 10652 17620 10658 17672
rect 11054 17620 11060 17672
rect 11112 17620 11118 17672
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17660 11299 17663
rect 11882 17660 11888 17672
rect 11287 17632 11888 17660
rect 11287 17629 11299 17632
rect 11241 17623 11299 17629
rect 11882 17620 11888 17632
rect 11940 17660 11946 17672
rect 12342 17660 12348 17672
rect 11940 17632 12348 17660
rect 11940 17620 11946 17632
rect 12342 17620 12348 17632
rect 12400 17620 12406 17672
rect 10612 17592 10640 17620
rect 10152 17564 10640 17592
rect 7432 17496 9260 17524
rect 9309 17527 9367 17533
rect 7432 17484 7438 17496
rect 9309 17493 9321 17527
rect 9355 17524 9367 17527
rect 9582 17524 9588 17536
rect 9355 17496 9588 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 11072 17524 11100 17620
rect 11701 17595 11759 17601
rect 11701 17561 11713 17595
rect 11747 17592 11759 17595
rect 12452 17592 12480 17768
rect 12526 17688 12532 17740
rect 12584 17688 12590 17740
rect 12636 17669 12664 17768
rect 16025 17765 16037 17768
rect 16071 17765 16083 17799
rect 16025 17759 16083 17765
rect 13354 17728 13360 17740
rect 13096 17700 13360 17728
rect 12621 17663 12679 17669
rect 12621 17629 12633 17663
rect 12667 17629 12679 17663
rect 12621 17623 12679 17629
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17629 12771 17663
rect 12713 17623 12771 17629
rect 12897 17663 12955 17669
rect 12897 17629 12909 17663
rect 12943 17629 12955 17663
rect 12897 17623 12955 17629
rect 12997 17663 13055 17669
rect 12997 17629 13009 17663
rect 13043 17660 13055 17663
rect 13096 17660 13124 17700
rect 13354 17688 13360 17700
rect 13412 17688 13418 17740
rect 13740 17700 14504 17728
rect 13740 17669 13768 17700
rect 14476 17672 14504 17700
rect 14642 17688 14648 17740
rect 14700 17688 14706 17740
rect 15102 17688 15108 17740
rect 15160 17728 15166 17740
rect 15473 17731 15531 17737
rect 15160 17700 15424 17728
rect 15160 17688 15166 17700
rect 13043 17632 13124 17660
rect 13173 17663 13231 17669
rect 13043 17629 13055 17632
rect 12997 17623 13055 17629
rect 13173 17629 13185 17663
rect 13219 17629 13231 17663
rect 13173 17623 13231 17629
rect 13725 17663 13783 17669
rect 13725 17629 13737 17663
rect 13771 17629 13783 17663
rect 13725 17623 13783 17629
rect 13909 17663 13967 17669
rect 13909 17629 13921 17663
rect 13955 17660 13967 17663
rect 14182 17660 14188 17672
rect 13955 17632 14188 17660
rect 13955 17629 13967 17632
rect 13909 17623 13967 17629
rect 11747 17564 12480 17592
rect 12728 17592 12756 17623
rect 12802 17592 12808 17604
rect 12728 17564 12808 17592
rect 11747 17561 11759 17564
rect 11701 17555 11759 17561
rect 12802 17552 12808 17564
rect 12860 17552 12866 17604
rect 12912 17592 12940 17623
rect 13188 17592 13216 17623
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 14277 17663 14335 17669
rect 14277 17629 14289 17663
rect 14323 17660 14335 17663
rect 14323 17632 14412 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 12912 17564 14044 17592
rect 14016 17536 14044 17564
rect 12158 17524 12164 17536
rect 11072 17496 12164 17524
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 12250 17484 12256 17536
rect 12308 17484 12314 17536
rect 12342 17484 12348 17536
rect 12400 17524 12406 17536
rect 12989 17527 13047 17533
rect 12989 17524 13001 17527
rect 12400 17496 13001 17524
rect 12400 17484 12406 17496
rect 12989 17493 13001 17496
rect 13035 17493 13047 17527
rect 12989 17487 13047 17493
rect 13078 17484 13084 17536
rect 13136 17524 13142 17536
rect 13630 17524 13636 17536
rect 13136 17496 13636 17524
rect 13136 17484 13142 17496
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 13998 17484 14004 17536
rect 14056 17484 14062 17536
rect 14200 17524 14228 17620
rect 14384 17604 14412 17632
rect 14458 17620 14464 17672
rect 14516 17620 14522 17672
rect 15396 17660 15424 17700
rect 15473 17697 15485 17731
rect 15519 17728 15531 17731
rect 15746 17728 15752 17740
rect 15519 17700 15752 17728
rect 15519 17697 15531 17700
rect 15473 17691 15531 17697
rect 15746 17688 15752 17700
rect 15804 17688 15810 17740
rect 16500 17728 16528 17836
rect 20625 17833 20637 17836
rect 20671 17864 20683 17867
rect 20806 17864 20812 17876
rect 20671 17836 20812 17864
rect 20671 17833 20683 17836
rect 20625 17827 20683 17833
rect 20806 17824 20812 17836
rect 20864 17864 20870 17876
rect 21634 17864 21640 17876
rect 20864 17836 21640 17864
rect 20864 17824 20870 17836
rect 21634 17824 21640 17836
rect 21692 17824 21698 17876
rect 22738 17824 22744 17876
rect 22796 17864 22802 17876
rect 22925 17867 22983 17873
rect 22925 17864 22937 17867
rect 22796 17836 22937 17864
rect 22796 17824 22802 17836
rect 22925 17833 22937 17836
rect 22971 17833 22983 17867
rect 22925 17827 22983 17833
rect 23290 17824 23296 17876
rect 23348 17864 23354 17876
rect 26878 17864 26884 17876
rect 23348 17836 26884 17864
rect 23348 17824 23354 17836
rect 26878 17824 26884 17836
rect 26936 17864 26942 17876
rect 27341 17867 27399 17873
rect 26936 17836 27108 17864
rect 26936 17824 26942 17836
rect 17218 17756 17224 17808
rect 17276 17796 17282 17808
rect 23658 17796 23664 17808
rect 17276 17768 23664 17796
rect 17276 17756 17282 17768
rect 23658 17756 23664 17768
rect 23716 17756 23722 17808
rect 23937 17799 23995 17805
rect 23937 17765 23949 17799
rect 23983 17796 23995 17799
rect 25593 17799 25651 17805
rect 23983 17768 25268 17796
rect 23983 17765 23995 17768
rect 23937 17759 23995 17765
rect 16408 17700 16528 17728
rect 15565 17663 15623 17669
rect 15565 17660 15577 17663
rect 14568 17632 15148 17660
rect 15396 17632 15577 17660
rect 14366 17552 14372 17604
rect 14424 17592 14430 17604
rect 14568 17592 14596 17632
rect 14424 17564 14596 17592
rect 15120 17592 15148 17632
rect 15565 17629 15577 17632
rect 15611 17629 15623 17663
rect 15565 17623 15623 17629
rect 15838 17620 15844 17672
rect 15896 17620 15902 17672
rect 16114 17620 16120 17672
rect 16172 17660 16178 17672
rect 16408 17669 16436 17700
rect 16574 17688 16580 17740
rect 16632 17728 16638 17740
rect 16632 17700 22508 17728
rect 16632 17688 16638 17700
rect 16255 17663 16313 17669
rect 16255 17660 16267 17663
rect 16172 17632 16267 17660
rect 16172 17620 16178 17632
rect 16255 17629 16267 17632
rect 16301 17629 16313 17663
rect 16255 17623 16313 17629
rect 16393 17663 16451 17669
rect 16393 17629 16405 17663
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 16485 17663 16543 17669
rect 16485 17629 16497 17663
rect 16531 17629 16543 17663
rect 16485 17623 16543 17629
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17660 16727 17663
rect 16758 17660 16764 17672
rect 16715 17632 16764 17660
rect 16715 17629 16727 17632
rect 16669 17623 16727 17629
rect 15378 17592 15384 17604
rect 15120 17564 15384 17592
rect 14424 17552 14430 17564
rect 15378 17552 15384 17564
rect 15436 17552 15442 17604
rect 15746 17552 15752 17604
rect 15804 17592 15810 17604
rect 15933 17595 15991 17601
rect 15933 17592 15945 17595
rect 15804 17564 15945 17592
rect 15804 17552 15810 17564
rect 15933 17561 15945 17564
rect 15979 17561 15991 17595
rect 15933 17555 15991 17561
rect 16408 17524 16436 17623
rect 14200 17496 16436 17524
rect 16500 17524 16528 17623
rect 16758 17620 16764 17632
rect 16816 17620 16822 17672
rect 16942 17620 16948 17672
rect 17000 17660 17006 17672
rect 17405 17663 17463 17669
rect 17405 17660 17417 17663
rect 17000 17632 17417 17660
rect 17000 17620 17006 17632
rect 17405 17629 17417 17632
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 17678 17620 17684 17672
rect 17736 17620 17742 17672
rect 17865 17663 17923 17669
rect 17865 17629 17877 17663
rect 17911 17629 17923 17663
rect 17865 17623 17923 17629
rect 17034 17552 17040 17604
rect 17092 17592 17098 17604
rect 17770 17592 17776 17604
rect 17092 17564 17776 17592
rect 17092 17552 17098 17564
rect 17770 17552 17776 17564
rect 17828 17592 17834 17604
rect 17880 17592 17908 17623
rect 18046 17620 18052 17672
rect 18104 17620 18110 17672
rect 18138 17620 18144 17672
rect 18196 17620 18202 17672
rect 18230 17620 18236 17672
rect 18288 17620 18294 17672
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17660 18475 17663
rect 18598 17660 18604 17672
rect 18463 17632 18604 17660
rect 18463 17629 18475 17632
rect 18417 17623 18475 17629
rect 18598 17620 18604 17632
rect 18656 17620 18662 17672
rect 18690 17620 18696 17672
rect 18748 17620 18754 17672
rect 18782 17620 18788 17672
rect 18840 17620 18846 17672
rect 18969 17663 19027 17669
rect 18969 17629 18981 17663
rect 19015 17660 19027 17663
rect 19334 17660 19340 17672
rect 19015 17632 19340 17660
rect 19015 17629 19027 17632
rect 18969 17623 19027 17629
rect 19334 17620 19340 17632
rect 19392 17620 19398 17672
rect 19426 17620 19432 17672
rect 19484 17660 19490 17672
rect 19978 17660 19984 17672
rect 19484 17632 19984 17660
rect 19484 17620 19490 17632
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 20162 17620 20168 17672
rect 20220 17660 20226 17672
rect 20349 17663 20407 17669
rect 20349 17660 20361 17663
rect 20220 17632 20361 17660
rect 20220 17620 20226 17632
rect 20349 17629 20361 17632
rect 20395 17660 20407 17663
rect 21174 17660 21180 17672
rect 20395 17632 21180 17660
rect 20395 17629 20407 17632
rect 20349 17623 20407 17629
rect 21174 17620 21180 17632
rect 21232 17620 21238 17672
rect 22094 17620 22100 17672
rect 22152 17620 22158 17672
rect 22278 17620 22284 17672
rect 22336 17620 22342 17672
rect 22480 17669 22508 17700
rect 23474 17688 23480 17740
rect 23532 17688 23538 17740
rect 24670 17688 24676 17740
rect 24728 17688 24734 17740
rect 24949 17731 25007 17737
rect 24949 17697 24961 17731
rect 24995 17728 25007 17731
rect 25133 17731 25191 17737
rect 25133 17728 25145 17731
rect 24995 17700 25145 17728
rect 24995 17697 25007 17700
rect 24949 17691 25007 17697
rect 25133 17697 25145 17700
rect 25179 17697 25191 17731
rect 25133 17691 25191 17697
rect 22465 17663 22523 17669
rect 22465 17629 22477 17663
rect 22511 17629 22523 17663
rect 22465 17623 22523 17629
rect 22557 17663 22615 17669
rect 22557 17629 22569 17663
rect 22603 17629 22615 17663
rect 22557 17623 22615 17629
rect 22649 17663 22707 17669
rect 22649 17629 22661 17663
rect 22695 17629 22707 17663
rect 22649 17623 22707 17629
rect 23569 17663 23627 17669
rect 23569 17629 23581 17663
rect 23615 17660 23627 17663
rect 24026 17660 24032 17672
rect 23615 17632 24032 17660
rect 23615 17629 23627 17632
rect 23569 17623 23627 17629
rect 18708 17592 18736 17620
rect 17828 17564 17908 17592
rect 18524 17564 18736 17592
rect 19996 17592 20024 17620
rect 20533 17595 20591 17601
rect 20533 17592 20545 17595
rect 19996 17564 20545 17592
rect 17828 17552 17834 17564
rect 17310 17524 17316 17536
rect 16500 17496 17316 17524
rect 17310 17484 17316 17496
rect 17368 17484 17374 17536
rect 17497 17527 17555 17533
rect 17497 17493 17509 17527
rect 17543 17524 17555 17527
rect 18524 17524 18552 17564
rect 20533 17561 20545 17564
rect 20579 17592 20591 17595
rect 20622 17592 20628 17604
rect 20579 17564 20628 17592
rect 20579 17561 20591 17564
rect 20533 17555 20591 17561
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 22112 17592 22140 17620
rect 22572 17592 22600 17623
rect 22112 17564 22600 17592
rect 22664 17592 22692 17623
rect 24026 17620 24032 17632
rect 24084 17620 24090 17672
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 24762 17660 24768 17672
rect 24627 17632 24768 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 24596 17592 24624 17623
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25240 17669 25268 17768
rect 25593 17765 25605 17799
rect 25639 17765 25651 17799
rect 25593 17759 25651 17765
rect 25225 17663 25283 17669
rect 25225 17629 25237 17663
rect 25271 17629 25283 17663
rect 25608 17660 25636 17759
rect 26234 17756 26240 17808
rect 26292 17756 26298 17808
rect 26605 17799 26663 17805
rect 26605 17765 26617 17799
rect 26651 17796 26663 17799
rect 27080 17796 27108 17836
rect 27341 17833 27353 17867
rect 27387 17864 27399 17867
rect 27982 17864 27988 17876
rect 27387 17836 27988 17864
rect 27387 17833 27399 17836
rect 27341 17827 27399 17833
rect 27982 17824 27988 17836
rect 28040 17824 28046 17876
rect 31202 17864 31208 17876
rect 28092 17836 31208 17864
rect 28092 17796 28120 17836
rect 31202 17824 31208 17836
rect 31260 17824 31266 17876
rect 31297 17867 31355 17873
rect 31297 17833 31309 17867
rect 31343 17864 31355 17867
rect 31386 17864 31392 17876
rect 31343 17836 31392 17864
rect 31343 17833 31355 17836
rect 31297 17827 31355 17833
rect 31386 17824 31392 17836
rect 31444 17824 31450 17876
rect 32125 17867 32183 17873
rect 32125 17833 32137 17867
rect 32171 17864 32183 17867
rect 32490 17864 32496 17876
rect 32171 17836 32496 17864
rect 32171 17833 32183 17836
rect 32125 17827 32183 17833
rect 32490 17824 32496 17836
rect 32548 17824 32554 17876
rect 29822 17796 29828 17808
rect 26651 17768 27016 17796
rect 27080 17768 28120 17796
rect 28184 17768 29828 17796
rect 26651 17765 26663 17768
rect 26605 17759 26663 17765
rect 26252 17728 26280 17756
rect 26988 17737 27016 17768
rect 26329 17731 26387 17737
rect 26329 17728 26341 17731
rect 26252 17700 26341 17728
rect 26329 17697 26341 17700
rect 26375 17697 26387 17731
rect 26329 17691 26387 17697
rect 26973 17731 27031 17737
rect 26973 17697 26985 17731
rect 27019 17697 27031 17731
rect 26973 17691 27031 17697
rect 27706 17688 27712 17740
rect 27764 17688 27770 17740
rect 28184 17728 28212 17768
rect 29822 17756 29828 17768
rect 29880 17796 29886 17808
rect 29880 17768 30236 17796
rect 29880 17756 29886 17768
rect 27816 17700 28212 17728
rect 27816 17672 27844 17700
rect 28258 17688 28264 17740
rect 28316 17728 28322 17740
rect 28316 17700 29960 17728
rect 28316 17688 28322 17700
rect 26237 17663 26295 17669
rect 26237 17660 26249 17663
rect 25608 17632 26249 17660
rect 25225 17623 25283 17629
rect 26237 17629 26249 17632
rect 26283 17629 26295 17663
rect 26237 17623 26295 17629
rect 27065 17663 27123 17669
rect 27065 17629 27077 17663
rect 27111 17629 27123 17663
rect 27065 17623 27123 17629
rect 22664 17564 24624 17592
rect 27080 17592 27108 17623
rect 27798 17620 27804 17672
rect 27856 17620 27862 17672
rect 27890 17620 27896 17672
rect 27948 17620 27954 17672
rect 27982 17620 27988 17672
rect 28040 17620 28046 17672
rect 28350 17620 28356 17672
rect 28408 17620 28414 17672
rect 28537 17663 28595 17669
rect 28537 17629 28549 17663
rect 28583 17629 28595 17663
rect 28537 17623 28595 17629
rect 27338 17592 27344 17604
rect 27080 17564 27344 17592
rect 27338 17552 27344 17564
rect 27396 17592 27402 17604
rect 28000 17592 28028 17620
rect 27396 17564 28028 17592
rect 27396 17552 27402 17564
rect 28166 17552 28172 17604
rect 28224 17592 28230 17604
rect 28552 17592 28580 17623
rect 28626 17620 28632 17672
rect 28684 17660 28690 17672
rect 29181 17663 29239 17669
rect 29181 17660 29193 17663
rect 28684 17632 29193 17660
rect 28684 17620 28690 17632
rect 29181 17629 29193 17632
rect 29227 17660 29239 17663
rect 29549 17663 29607 17669
rect 29549 17660 29561 17663
rect 29227 17632 29561 17660
rect 29227 17629 29239 17632
rect 29181 17623 29239 17629
rect 29549 17629 29561 17632
rect 29595 17629 29607 17663
rect 29549 17623 29607 17629
rect 29730 17620 29736 17672
rect 29788 17620 29794 17672
rect 29932 17669 29960 17700
rect 29825 17663 29883 17669
rect 29825 17629 29837 17663
rect 29871 17629 29883 17663
rect 29825 17623 29883 17629
rect 29917 17663 29975 17669
rect 29917 17629 29929 17663
rect 29963 17660 29975 17663
rect 30098 17660 30104 17672
rect 29963 17632 30104 17660
rect 29963 17629 29975 17632
rect 29917 17623 29975 17629
rect 28224 17564 28580 17592
rect 29840 17592 29868 17623
rect 30098 17620 30104 17632
rect 30156 17620 30162 17672
rect 30208 17660 30236 17768
rect 30282 17756 30288 17808
rect 30340 17796 30346 17808
rect 32582 17796 32588 17808
rect 30340 17768 32588 17796
rect 30340 17756 30346 17768
rect 30282 17660 30288 17672
rect 30208 17632 30288 17660
rect 30282 17620 30288 17632
rect 30340 17620 30346 17672
rect 30484 17669 30512 17768
rect 32582 17756 32588 17768
rect 32640 17756 32646 17808
rect 34054 17756 34060 17808
rect 34112 17756 34118 17808
rect 31294 17688 31300 17740
rect 31352 17688 31358 17740
rect 30469 17663 30527 17669
rect 30469 17629 30481 17663
rect 30515 17629 30527 17663
rect 30469 17623 30527 17629
rect 31205 17663 31263 17669
rect 31205 17629 31217 17663
rect 31251 17660 31263 17663
rect 31312 17660 31340 17688
rect 31251 17632 31340 17660
rect 31251 17629 31263 17632
rect 31205 17623 31263 17629
rect 32030 17620 32036 17672
rect 32088 17620 32094 17672
rect 33410 17620 33416 17672
rect 33468 17660 33474 17672
rect 33781 17663 33839 17669
rect 33781 17660 33793 17663
rect 33468 17632 33793 17660
rect 33468 17620 33474 17632
rect 33781 17629 33793 17632
rect 33827 17629 33839 17663
rect 33781 17623 33839 17629
rect 33962 17620 33968 17672
rect 34020 17660 34026 17672
rect 34057 17663 34115 17669
rect 34057 17660 34069 17663
rect 34020 17632 34069 17660
rect 34020 17620 34026 17632
rect 34057 17629 34069 17632
rect 34103 17629 34115 17663
rect 34057 17623 34115 17629
rect 29840 17564 30420 17592
rect 28224 17552 28230 17564
rect 17543 17496 18552 17524
rect 17543 17493 17555 17496
rect 17497 17487 17555 17493
rect 18598 17484 18604 17536
rect 18656 17484 18662 17536
rect 18874 17484 18880 17536
rect 18932 17484 18938 17536
rect 18966 17484 18972 17536
rect 19024 17524 19030 17536
rect 29178 17524 29184 17536
rect 19024 17496 29184 17524
rect 19024 17484 19030 17496
rect 29178 17484 29184 17496
rect 29236 17484 29242 17536
rect 30190 17484 30196 17536
rect 30248 17484 30254 17536
rect 30392 17533 30420 17564
rect 30377 17527 30435 17533
rect 30377 17493 30389 17527
rect 30423 17524 30435 17527
rect 31846 17524 31852 17536
rect 30423 17496 31852 17524
rect 30423 17493 30435 17496
rect 30377 17487 30435 17493
rect 31846 17484 31852 17496
rect 31904 17484 31910 17536
rect 33778 17484 33784 17536
rect 33836 17524 33842 17536
rect 33873 17527 33931 17533
rect 33873 17524 33885 17527
rect 33836 17496 33885 17524
rect 33836 17484 33842 17496
rect 33873 17493 33885 17496
rect 33919 17493 33931 17527
rect 33873 17487 33931 17493
rect 1104 17434 38272 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38272 17434
rect 1104 17360 38272 17382
rect 3418 17280 3424 17332
rect 3476 17280 3482 17332
rect 4246 17280 4252 17332
rect 4304 17280 4310 17332
rect 4525 17323 4583 17329
rect 4525 17289 4537 17323
rect 4571 17289 4583 17323
rect 4525 17283 4583 17289
rect 4062 17212 4068 17264
rect 4120 17212 4126 17264
rect 3053 17187 3111 17193
rect 3053 17153 3065 17187
rect 3099 17153 3111 17187
rect 3053 17147 3111 17153
rect 3068 17116 3096 17147
rect 3234 17144 3240 17196
rect 3292 17144 3298 17196
rect 3786 17116 3792 17128
rect 3068 17088 3792 17116
rect 3786 17076 3792 17088
rect 3844 17116 3850 17128
rect 4080 17116 4108 17212
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 4540 17184 4568 17283
rect 5718 17280 5724 17332
rect 5776 17280 5782 17332
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 6549 17323 6607 17329
rect 6549 17320 6561 17323
rect 6420 17292 6561 17320
rect 6420 17280 6426 17292
rect 6549 17289 6561 17292
rect 6595 17289 6607 17323
rect 6549 17283 6607 17289
rect 6917 17323 6975 17329
rect 6917 17289 6929 17323
rect 6963 17289 6975 17323
rect 6917 17283 6975 17289
rect 7377 17323 7435 17329
rect 7377 17289 7389 17323
rect 7423 17320 7435 17323
rect 7742 17320 7748 17332
rect 7423 17292 7748 17320
rect 7423 17289 7435 17292
rect 7377 17283 7435 17289
rect 4798 17212 4804 17264
rect 4856 17252 4862 17264
rect 4893 17255 4951 17261
rect 4893 17252 4905 17255
rect 4856 17224 4905 17252
rect 4856 17212 4862 17224
rect 4893 17221 4905 17224
rect 4939 17252 4951 17255
rect 5736 17252 5764 17280
rect 5905 17255 5963 17261
rect 5905 17252 5917 17255
rect 4939 17224 5917 17252
rect 4939 17221 4951 17224
rect 4893 17215 4951 17221
rect 5905 17221 5917 17224
rect 5951 17221 5963 17255
rect 5905 17215 5963 17221
rect 5721 17187 5779 17193
rect 5721 17184 5733 17187
rect 4479 17156 4568 17184
rect 4908 17156 5733 17184
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 4908 17116 4936 17156
rect 5721 17153 5733 17156
rect 5767 17153 5779 17187
rect 5721 17147 5779 17153
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 6932 17184 6960 17283
rect 7742 17280 7748 17292
rect 7800 17280 7806 17332
rect 9490 17320 9496 17332
rect 8956 17292 9496 17320
rect 6779 17156 6960 17184
rect 7285 17187 7343 17193
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 8478 17184 8484 17196
rect 7331 17156 8484 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 8478 17144 8484 17156
rect 8536 17144 8542 17196
rect 8956 17193 8984 17292
rect 9490 17280 9496 17292
rect 9548 17320 9554 17332
rect 10134 17320 10140 17332
rect 9548 17292 10140 17320
rect 9548 17280 9554 17292
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 11146 17320 11152 17332
rect 10244 17292 11152 17320
rect 9398 17212 9404 17264
rect 9456 17212 9462 17264
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 9953 17255 10011 17261
rect 9953 17252 9965 17255
rect 9732 17224 9965 17252
rect 9732 17212 9738 17224
rect 9953 17221 9965 17224
rect 9999 17221 10011 17255
rect 9953 17215 10011 17221
rect 10244 17215 10272 17292
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 11974 17280 11980 17332
rect 12032 17280 12038 17332
rect 12250 17320 12256 17332
rect 12084 17292 12256 17320
rect 8941 17187 8999 17193
rect 8941 17153 8953 17187
rect 8987 17153 8999 17187
rect 8941 17147 8999 17153
rect 9125 17187 9183 17193
rect 9125 17153 9137 17187
rect 9171 17184 9183 17187
rect 9416 17184 9444 17212
rect 9171 17156 9444 17184
rect 10228 17209 10286 17215
rect 10318 17212 10324 17264
rect 10376 17212 10382 17264
rect 12084 17252 12112 17292
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 12434 17280 12440 17332
rect 12492 17280 12498 17332
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 15562 17320 15568 17332
rect 14056 17292 15568 17320
rect 14056 17280 14062 17292
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 16206 17280 16212 17332
rect 16264 17320 16270 17332
rect 16758 17320 16764 17332
rect 16264 17292 16764 17320
rect 16264 17280 16270 17292
rect 16758 17280 16764 17292
rect 16816 17320 16822 17332
rect 16816 17292 18736 17320
rect 16816 17280 16822 17292
rect 12452 17252 12480 17280
rect 17218 17252 17224 17264
rect 10980 17224 12112 17252
rect 12176 17224 12480 17252
rect 13924 17224 17224 17252
rect 10228 17175 10240 17209
rect 10274 17175 10286 17209
rect 10228 17169 10286 17175
rect 10320 17209 10378 17212
rect 10320 17175 10332 17209
rect 10366 17175 10378 17209
rect 10320 17169 10378 17175
rect 9171 17153 9183 17156
rect 9125 17147 9183 17153
rect 10410 17144 10416 17196
rect 10468 17144 10474 17196
rect 10594 17144 10600 17196
rect 10652 17184 10658 17196
rect 10980 17184 11008 17224
rect 10652 17156 11008 17184
rect 10652 17144 10658 17156
rect 11606 17144 11612 17196
rect 11664 17144 11670 17196
rect 11790 17144 11796 17196
rect 11848 17184 11854 17196
rect 12176 17193 12204 17224
rect 11977 17187 12035 17193
rect 11977 17184 11989 17187
rect 11848 17156 11989 17184
rect 11848 17144 11854 17156
rect 11977 17153 11989 17156
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 12250 17144 12256 17196
rect 12308 17144 12314 17196
rect 12437 17187 12495 17193
rect 12437 17153 12449 17187
rect 12483 17184 12495 17187
rect 12618 17184 12624 17196
rect 12483 17156 12624 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 3844 17088 4936 17116
rect 3844 17076 3850 17088
rect 4982 17076 4988 17128
rect 5040 17076 5046 17128
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17085 5135 17119
rect 5077 17079 5135 17085
rect 3050 17008 3056 17060
rect 3108 17048 3114 17060
rect 5092 17048 5120 17079
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7469 17119 7527 17125
rect 7469 17116 7481 17119
rect 7248 17088 7481 17116
rect 7248 17076 7254 17088
rect 7469 17085 7481 17088
rect 7515 17085 7527 17119
rect 11624 17116 11652 17144
rect 12342 17116 12348 17128
rect 11624 17088 12348 17116
rect 7469 17079 7527 17085
rect 12342 17076 12348 17088
rect 12400 17076 12406 17128
rect 3108 17020 5120 17048
rect 3108 17008 3114 17020
rect 7558 17008 7564 17060
rect 7616 17048 7622 17060
rect 13924 17048 13952 17224
rect 17218 17212 17224 17224
rect 17276 17212 17282 17264
rect 18708 17252 18736 17292
rect 19058 17280 19064 17332
rect 19116 17320 19122 17332
rect 19426 17320 19432 17332
rect 19116 17292 19432 17320
rect 19116 17280 19122 17292
rect 19426 17280 19432 17292
rect 19484 17320 19490 17332
rect 19702 17320 19708 17332
rect 19484 17292 19708 17320
rect 19484 17280 19490 17292
rect 19702 17280 19708 17292
rect 19760 17280 19766 17332
rect 21082 17320 21088 17332
rect 19904 17292 21088 17320
rect 19904 17261 19932 17292
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 23290 17320 23296 17332
rect 22388 17292 23296 17320
rect 19889 17255 19947 17261
rect 19889 17252 19901 17255
rect 18708 17224 19901 17252
rect 19889 17221 19901 17224
rect 19935 17221 19947 17255
rect 19889 17215 19947 17221
rect 19978 17212 19984 17264
rect 20036 17212 20042 17264
rect 20162 17252 20168 17264
rect 20093 17224 20168 17252
rect 15562 17144 15568 17196
rect 15620 17184 15626 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 15620 17156 16681 17184
rect 15620 17144 15626 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17184 16911 17187
rect 17862 17184 17868 17196
rect 16899 17156 17868 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 17862 17144 17868 17156
rect 17920 17184 17926 17196
rect 18322 17184 18328 17196
rect 17920 17156 18328 17184
rect 17920 17144 17926 17156
rect 18322 17144 18328 17156
rect 18380 17144 18386 17196
rect 18966 17144 18972 17196
rect 19024 17144 19030 17196
rect 19610 17144 19616 17196
rect 19668 17144 19674 17196
rect 19702 17144 19708 17196
rect 19760 17184 19766 17196
rect 20093 17193 20121 17224
rect 20162 17212 20168 17224
rect 20220 17212 20226 17264
rect 20346 17212 20352 17264
rect 20404 17212 20410 17264
rect 20078 17187 20136 17193
rect 20078 17184 20090 17187
rect 19760 17156 19805 17184
rect 20036 17156 20090 17184
rect 19760 17144 19766 17156
rect 20078 17153 20090 17156
rect 20124 17153 20136 17187
rect 20625 17187 20683 17193
rect 20625 17184 20637 17187
rect 20078 17147 20136 17153
rect 20180 17156 20637 17184
rect 14461 17119 14519 17125
rect 14461 17085 14473 17119
rect 14507 17116 14519 17119
rect 14550 17116 14556 17128
rect 14507 17088 14556 17116
rect 14507 17085 14519 17088
rect 14461 17079 14519 17085
rect 14550 17076 14556 17088
rect 14608 17076 14614 17128
rect 15746 17076 15752 17128
rect 15804 17116 15810 17128
rect 16942 17116 16948 17128
rect 15804 17088 16948 17116
rect 15804 17076 15810 17088
rect 16942 17076 16948 17088
rect 17000 17076 17006 17128
rect 7616 17020 13952 17048
rect 14185 17051 14243 17057
rect 7616 17008 7622 17020
rect 14185 17017 14197 17051
rect 14231 17048 14243 17051
rect 14366 17048 14372 17060
rect 14231 17020 14372 17048
rect 14231 17017 14243 17020
rect 14185 17011 14243 17017
rect 14366 17008 14372 17020
rect 14424 17008 14430 17060
rect 18984 17048 19012 17144
rect 20093 17116 20121 17147
rect 20180 17128 20208 17156
rect 20625 17153 20637 17156
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17153 20775 17187
rect 20717 17147 20775 17153
rect 16592 17020 19012 17048
rect 19306 17088 20121 17116
rect 6086 16940 6092 16992
rect 6144 16940 6150 16992
rect 9309 16983 9367 16989
rect 9309 16949 9321 16983
rect 9355 16980 9367 16983
rect 9582 16980 9588 16992
rect 9355 16952 9588 16980
rect 9355 16949 9367 16952
rect 9309 16943 9367 16949
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 11790 16940 11796 16992
rect 11848 16980 11854 16992
rect 16592 16980 16620 17020
rect 11848 16952 16620 16980
rect 11848 16940 11854 16952
rect 16666 16940 16672 16992
rect 16724 16940 16730 16992
rect 17037 16983 17095 16989
rect 17037 16949 17049 16983
rect 17083 16980 17095 16983
rect 18230 16980 18236 16992
rect 17083 16952 18236 16980
rect 17083 16949 17095 16952
rect 17037 16943 17095 16949
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 18690 16940 18696 16992
rect 18748 16980 18754 16992
rect 19306 16980 19334 17088
rect 20162 17076 20168 17128
rect 20220 17076 20226 17128
rect 20530 17076 20536 17128
rect 20588 17116 20594 17128
rect 20732 17116 20760 17147
rect 20806 17144 20812 17196
rect 20864 17193 20870 17196
rect 22388 17193 22416 17292
rect 23290 17280 23296 17292
rect 23348 17280 23354 17332
rect 23474 17280 23480 17332
rect 23532 17280 23538 17332
rect 28350 17280 28356 17332
rect 28408 17280 28414 17332
rect 28460 17292 28672 17320
rect 23492 17252 23520 17280
rect 28261 17255 28319 17261
rect 22756 17224 23520 17252
rect 28000 17224 28205 17252
rect 20864 17184 20872 17193
rect 20993 17187 21051 17193
rect 20864 17156 20909 17184
rect 20864 17147 20872 17156
rect 20993 17153 21005 17187
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 22373 17187 22431 17193
rect 22373 17153 22385 17187
rect 22419 17153 22431 17187
rect 22373 17147 22431 17153
rect 20864 17144 20870 17147
rect 20588 17088 20760 17116
rect 20588 17076 20594 17088
rect 20714 17048 20720 17060
rect 20180 17020 20720 17048
rect 18748 16952 19334 16980
rect 18748 16940 18754 16952
rect 19794 16940 19800 16992
rect 19852 16980 19858 16992
rect 20180 16980 20208 17020
rect 20714 17008 20720 17020
rect 20772 17008 20778 17060
rect 19852 16952 20208 16980
rect 20257 16983 20315 16989
rect 19852 16940 19858 16952
rect 20257 16949 20269 16983
rect 20303 16980 20315 16983
rect 21008 16980 21036 17147
rect 22756 17125 22784 17224
rect 22922 17144 22928 17196
rect 22980 17144 22986 17196
rect 23477 17187 23535 17193
rect 23477 17153 23489 17187
rect 23523 17184 23535 17187
rect 27798 17184 27804 17196
rect 23523 17156 27804 17184
rect 23523 17153 23535 17156
rect 23477 17147 23535 17153
rect 27798 17144 27804 17156
rect 27856 17144 27862 17196
rect 28000 17193 28028 17224
rect 27985 17187 28043 17193
rect 27985 17153 27997 17187
rect 28031 17153 28043 17187
rect 27985 17147 28043 17153
rect 28077 17187 28135 17193
rect 28077 17153 28089 17187
rect 28123 17153 28135 17187
rect 28177 17184 28205 17224
rect 28261 17221 28273 17255
rect 28307 17252 28319 17255
rect 28460 17252 28488 17292
rect 28644 17264 28672 17292
rect 29178 17280 29184 17332
rect 29236 17280 29242 17332
rect 30190 17280 30196 17332
rect 30248 17280 30254 17332
rect 32030 17320 32036 17332
rect 31680 17292 32036 17320
rect 28307 17224 28488 17252
rect 28521 17255 28579 17261
rect 28307 17221 28319 17224
rect 28261 17215 28319 17221
rect 28521 17221 28533 17255
rect 28567 17252 28579 17255
rect 28567 17221 28580 17252
rect 28521 17215 28580 17221
rect 28552 17184 28580 17215
rect 28626 17212 28632 17264
rect 28684 17252 28690 17264
rect 28721 17255 28779 17261
rect 28721 17252 28733 17255
rect 28684 17224 28733 17252
rect 28684 17212 28690 17224
rect 28721 17221 28733 17224
rect 28767 17221 28779 17255
rect 30208 17252 30236 17280
rect 31680 17261 31708 17292
rect 32030 17280 32036 17292
rect 32088 17320 32094 17332
rect 32088 17292 32536 17320
rect 32088 17280 32094 17292
rect 28721 17215 28779 17221
rect 29012 17224 30236 17252
rect 31665 17255 31723 17261
rect 29012 17193 29040 17224
rect 31665 17221 31677 17255
rect 31711 17221 31723 17255
rect 31665 17215 31723 17221
rect 32508 17218 32536 17292
rect 32858 17280 32864 17332
rect 32916 17320 32922 17332
rect 33042 17320 33048 17332
rect 32916 17292 33048 17320
rect 32916 17280 32922 17292
rect 33042 17280 33048 17292
rect 33100 17320 33106 17332
rect 33137 17323 33195 17329
rect 33137 17320 33149 17323
rect 33100 17292 33149 17320
rect 33100 17280 33106 17292
rect 33137 17289 33149 17292
rect 33183 17289 33195 17323
rect 33137 17283 33195 17289
rect 33962 17280 33968 17332
rect 34020 17329 34026 17332
rect 34020 17323 34039 17329
rect 34027 17289 34039 17323
rect 34020 17283 34039 17289
rect 34149 17323 34207 17329
rect 34149 17289 34161 17323
rect 34195 17289 34207 17323
rect 34149 17283 34207 17289
rect 34020 17280 34026 17283
rect 28177 17156 28580 17184
rect 28077 17147 28135 17153
rect 22465 17119 22523 17125
rect 22465 17085 22477 17119
rect 22511 17085 22523 17119
rect 22465 17079 22523 17085
rect 22741 17119 22799 17125
rect 22741 17085 22753 17119
rect 22787 17085 22799 17119
rect 22741 17079 22799 17085
rect 22480 17048 22508 17079
rect 23106 17076 23112 17128
rect 23164 17076 23170 17128
rect 28092 17116 28120 17147
rect 28552 17116 28580 17156
rect 28997 17187 29055 17193
rect 28997 17153 29009 17187
rect 29043 17153 29055 17187
rect 28997 17147 29055 17153
rect 29178 17144 29184 17196
rect 29236 17144 29242 17196
rect 29549 17187 29607 17193
rect 29549 17153 29561 17187
rect 29595 17184 29607 17187
rect 29638 17184 29644 17196
rect 29595 17156 29644 17184
rect 29595 17153 29607 17156
rect 29549 17147 29607 17153
rect 29638 17144 29644 17156
rect 29696 17144 29702 17196
rect 31846 17144 31852 17196
rect 31904 17144 31910 17196
rect 31941 17187 31999 17193
rect 31941 17153 31953 17187
rect 31987 17184 31999 17187
rect 32122 17184 32128 17196
rect 31987 17156 32128 17184
rect 31987 17153 31999 17156
rect 31941 17147 31999 17153
rect 32122 17144 32128 17156
rect 32180 17144 32186 17196
rect 32416 17193 32536 17218
rect 33778 17212 33784 17264
rect 33836 17212 33842 17264
rect 32400 17190 32536 17193
rect 32400 17187 32458 17190
rect 32400 17153 32412 17187
rect 32446 17153 32458 17187
rect 32400 17147 32458 17153
rect 32858 17144 32864 17196
rect 32916 17144 32922 17196
rect 33045 17187 33103 17193
rect 33045 17153 33057 17187
rect 33091 17153 33103 17187
rect 34164 17184 34192 17283
rect 34514 17212 34520 17264
rect 34572 17252 34578 17264
rect 34572 17224 35204 17252
rect 34572 17212 34578 17224
rect 34425 17187 34483 17193
rect 34425 17184 34437 17187
rect 34164 17156 34437 17184
rect 33045 17147 33103 17153
rect 34425 17153 34437 17156
rect 34471 17184 34483 17187
rect 34885 17187 34943 17193
rect 34471 17156 34652 17184
rect 34471 17153 34483 17156
rect 34425 17147 34483 17153
rect 28092 17088 28488 17116
rect 28552 17088 29408 17116
rect 23124 17048 23152 17076
rect 22480 17020 23152 17048
rect 23290 17008 23296 17060
rect 23348 17048 23354 17060
rect 25130 17048 25136 17060
rect 23348 17020 25136 17048
rect 23348 17008 23354 17020
rect 25130 17008 25136 17020
rect 25188 17008 25194 17060
rect 28166 17008 28172 17060
rect 28224 17048 28230 17060
rect 28261 17051 28319 17057
rect 28261 17048 28273 17051
rect 28224 17020 28273 17048
rect 28224 17008 28230 17020
rect 28261 17017 28273 17020
rect 28307 17017 28319 17051
rect 28261 17011 28319 17017
rect 20303 16952 21036 16980
rect 20303 16949 20315 16952
rect 20257 16943 20315 16949
rect 24578 16940 24584 16992
rect 24636 16980 24642 16992
rect 28074 16980 28080 16992
rect 24636 16952 28080 16980
rect 24636 16940 24642 16952
rect 28074 16940 28080 16952
rect 28132 16940 28138 16992
rect 28460 16980 28488 17088
rect 29380 16992 29408 17088
rect 30098 17076 30104 17128
rect 30156 17116 30162 17128
rect 30156 17108 32260 17116
rect 32306 17108 32312 17128
rect 30156 17088 32312 17108
rect 30156 17076 30162 17088
rect 32232 17080 32312 17088
rect 32306 17076 32312 17080
rect 32364 17076 32370 17128
rect 32493 17119 32551 17125
rect 32493 17108 32505 17119
rect 32416 17085 32505 17108
rect 32539 17085 32551 17119
rect 32416 17080 32551 17085
rect 31665 17051 31723 17057
rect 31665 17017 31677 17051
rect 31711 17048 31723 17051
rect 32030 17048 32036 17060
rect 31711 17020 32036 17048
rect 31711 17017 31723 17020
rect 31665 17011 31723 17017
rect 32030 17008 32036 17020
rect 32088 17008 32094 17060
rect 28537 16983 28595 16989
rect 28537 16980 28549 16983
rect 28460 16952 28549 16980
rect 28537 16949 28549 16952
rect 28583 16980 28595 16983
rect 29270 16980 29276 16992
rect 28583 16952 29276 16980
rect 28583 16949 28595 16952
rect 28537 16943 28595 16949
rect 29270 16940 29276 16952
rect 29328 16940 29334 16992
rect 29362 16940 29368 16992
rect 29420 16940 29426 16992
rect 30282 16940 30288 16992
rect 30340 16980 30346 16992
rect 31754 16980 31760 16992
rect 30340 16952 31760 16980
rect 30340 16940 30346 16952
rect 31754 16940 31760 16952
rect 31812 16940 31818 16992
rect 31846 16940 31852 16992
rect 31904 16980 31910 16992
rect 32416 16980 32444 17080
rect 32493 17079 32551 17080
rect 32582 17076 32588 17128
rect 32640 17076 32646 17128
rect 32769 17119 32827 17125
rect 32769 17085 32781 17119
rect 32815 17116 32827 17119
rect 33060 17116 33088 17147
rect 32815 17088 33088 17116
rect 32815 17085 32827 17088
rect 32769 17079 32827 17085
rect 34054 17076 34060 17128
rect 34112 17076 34118 17128
rect 34514 17076 34520 17128
rect 34572 17076 34578 17128
rect 34624 17116 34652 17156
rect 34885 17153 34897 17187
rect 34931 17184 34943 17187
rect 34931 17156 35112 17184
rect 34931 17153 34943 17156
rect 34885 17147 34943 17153
rect 34977 17119 35035 17125
rect 34977 17116 34989 17119
rect 34624 17088 34989 17116
rect 34977 17085 34989 17088
rect 35023 17085 35035 17119
rect 34977 17079 35035 17085
rect 31904 16952 32444 16980
rect 31904 16940 31910 16952
rect 33410 16940 33416 16992
rect 33468 16980 33474 16992
rect 33965 16983 34023 16989
rect 33965 16980 33977 16983
rect 33468 16952 33977 16980
rect 33468 16940 33474 16952
rect 33965 16949 33977 16952
rect 34011 16949 34023 16983
rect 34072 16980 34100 17076
rect 35084 17048 35112 17156
rect 35176 17125 35204 17224
rect 35161 17119 35219 17125
rect 35161 17085 35173 17119
rect 35207 17085 35219 17119
rect 35161 17079 35219 17085
rect 34440 17020 35112 17048
rect 34440 16989 34468 17020
rect 34425 16983 34483 16989
rect 34425 16980 34437 16983
rect 34072 16952 34437 16980
rect 33965 16943 34023 16949
rect 34425 16949 34437 16952
rect 34471 16949 34483 16983
rect 34425 16943 34483 16949
rect 34790 16940 34796 16992
rect 34848 16940 34854 16992
rect 35069 16983 35127 16989
rect 35069 16949 35081 16983
rect 35115 16980 35127 16983
rect 35342 16980 35348 16992
rect 35115 16952 35348 16980
rect 35115 16949 35127 16952
rect 35069 16943 35127 16949
rect 35342 16940 35348 16952
rect 35400 16940 35406 16992
rect 1104 16890 38272 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38272 16890
rect 1104 16816 38272 16838
rect 3602 16736 3608 16788
rect 3660 16776 3666 16788
rect 3660 16748 4660 16776
rect 3660 16736 3666 16748
rect 3789 16711 3847 16717
rect 3789 16708 3801 16711
rect 2792 16680 3801 16708
rect 2792 16649 2820 16680
rect 3789 16677 3801 16680
rect 3835 16677 3847 16711
rect 3789 16671 3847 16677
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16609 2835 16643
rect 2777 16603 2835 16609
rect 2961 16643 3019 16649
rect 2961 16609 2973 16643
rect 3007 16640 3019 16643
rect 3050 16640 3056 16652
rect 3007 16612 3056 16640
rect 3007 16609 3019 16612
rect 2961 16603 3019 16609
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 4430 16600 4436 16652
rect 4488 16600 4494 16652
rect 1949 16575 2007 16581
rect 1949 16541 1961 16575
rect 1995 16572 2007 16575
rect 2130 16572 2136 16584
rect 1995 16544 2136 16572
rect 1995 16541 2007 16544
rect 1949 16535 2007 16541
rect 2130 16532 2136 16544
rect 2188 16532 2194 16584
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16572 2283 16575
rect 2271 16544 2360 16572
rect 2271 16541 2283 16544
rect 2225 16535 2283 16541
rect 1762 16396 1768 16448
rect 1820 16396 1826 16448
rect 1946 16396 1952 16448
rect 2004 16436 2010 16448
rect 2332 16445 2360 16544
rect 3970 16532 3976 16584
rect 4028 16532 4034 16584
rect 4154 16532 4160 16584
rect 4212 16574 4218 16584
rect 4517 16575 4575 16581
rect 4212 16572 4384 16574
rect 4212 16546 4476 16572
rect 4212 16532 4218 16546
rect 4356 16544 4476 16546
rect 4065 16507 4123 16513
rect 4065 16473 4077 16507
rect 4111 16473 4123 16507
rect 4065 16467 4123 16473
rect 2041 16439 2099 16445
rect 2041 16436 2053 16439
rect 2004 16408 2053 16436
rect 2004 16396 2010 16408
rect 2041 16405 2053 16408
rect 2087 16405 2099 16439
rect 2041 16399 2099 16405
rect 2317 16439 2375 16445
rect 2317 16405 2329 16439
rect 2363 16405 2375 16439
rect 2317 16399 2375 16405
rect 2685 16439 2743 16445
rect 2685 16405 2697 16439
rect 2731 16436 2743 16439
rect 3142 16436 3148 16448
rect 2731 16408 3148 16436
rect 2731 16405 2743 16408
rect 2685 16399 2743 16405
rect 3142 16396 3148 16408
rect 3200 16396 3206 16448
rect 4080 16436 4108 16467
rect 4246 16464 4252 16516
rect 4304 16513 4310 16516
rect 4304 16507 4353 16513
rect 4304 16473 4307 16507
rect 4341 16473 4353 16507
rect 4448 16504 4476 16544
rect 4517 16541 4529 16575
rect 4563 16572 4575 16575
rect 4632 16572 4660 16748
rect 6086 16736 6092 16788
rect 6144 16776 6150 16788
rect 6144 16748 12434 16776
rect 6144 16736 6150 16748
rect 8389 16711 8447 16717
rect 8389 16677 8401 16711
rect 8435 16708 8447 16711
rect 8478 16708 8484 16720
rect 8435 16680 8484 16708
rect 8435 16677 8447 16680
rect 8389 16671 8447 16677
rect 8478 16668 8484 16680
rect 8536 16668 8542 16720
rect 8588 16680 9260 16708
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 8588 16640 8616 16680
rect 8352 16612 8616 16640
rect 8352 16600 8358 16612
rect 8588 16581 8616 16612
rect 8846 16600 8852 16652
rect 8904 16640 8910 16652
rect 9125 16643 9183 16649
rect 9125 16640 9137 16643
rect 8904 16612 9137 16640
rect 8904 16600 8910 16612
rect 9125 16609 9137 16612
rect 9171 16609 9183 16643
rect 9232 16640 9260 16680
rect 11974 16668 11980 16720
rect 12032 16708 12038 16720
rect 12250 16708 12256 16720
rect 12032 16680 12256 16708
rect 12032 16668 12038 16680
rect 12250 16668 12256 16680
rect 12308 16668 12314 16720
rect 12406 16708 12434 16748
rect 14274 16736 14280 16788
rect 14332 16776 14338 16788
rect 16485 16779 16543 16785
rect 16485 16776 16497 16779
rect 14332 16748 16497 16776
rect 14332 16736 14338 16748
rect 16485 16745 16497 16748
rect 16531 16745 16543 16779
rect 16485 16739 16543 16745
rect 16574 16736 16580 16788
rect 16632 16736 16638 16788
rect 16666 16736 16672 16788
rect 16724 16736 16730 16788
rect 19334 16776 19340 16788
rect 18248 16748 19340 16776
rect 16592 16708 16620 16736
rect 12406 16680 16620 16708
rect 9398 16640 9404 16652
rect 9232 16612 9404 16640
rect 9125 16603 9183 16609
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 15654 16600 15660 16652
rect 15712 16640 15718 16652
rect 16117 16643 16175 16649
rect 16117 16640 16129 16643
rect 15712 16612 16129 16640
rect 15712 16600 15718 16612
rect 16117 16609 16129 16612
rect 16163 16609 16175 16643
rect 16117 16603 16175 16609
rect 4563 16544 4660 16572
rect 8573 16575 8631 16581
rect 4563 16541 4575 16544
rect 4517 16535 4575 16541
rect 8573 16541 8585 16575
rect 8619 16541 8631 16575
rect 8573 16535 8631 16541
rect 8757 16575 8815 16581
rect 8757 16541 8769 16575
rect 8803 16572 8815 16575
rect 8938 16572 8944 16584
rect 8803 16544 8944 16572
rect 8803 16541 8815 16544
rect 8757 16535 8815 16541
rect 8938 16532 8944 16544
rect 8996 16532 9002 16584
rect 14550 16532 14556 16584
rect 14608 16572 14614 16584
rect 14737 16575 14795 16581
rect 14737 16572 14749 16575
rect 14608 16544 14749 16572
rect 14608 16532 14614 16544
rect 14737 16541 14749 16544
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 15378 16532 15384 16584
rect 15436 16532 15442 16584
rect 15838 16532 15844 16584
rect 15896 16532 15902 16584
rect 16684 16572 16712 16736
rect 17494 16708 17500 16720
rect 17236 16680 17500 16708
rect 16850 16572 16856 16584
rect 16684 16544 16856 16572
rect 16850 16532 16856 16544
rect 16908 16572 16914 16584
rect 17236 16581 17264 16680
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 17310 16600 17316 16652
rect 17368 16640 17374 16652
rect 17368 16612 17908 16640
rect 17368 16600 17374 16612
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16908 16544 16957 16572
rect 16908 16532 16914 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 16945 16535 17003 16541
rect 17221 16575 17279 16581
rect 17221 16541 17233 16575
rect 17267 16541 17279 16575
rect 17221 16535 17279 16541
rect 17586 16532 17592 16584
rect 17644 16532 17650 16584
rect 5902 16504 5908 16516
rect 4448 16476 5908 16504
rect 4304 16467 4353 16473
rect 4304 16464 4310 16467
rect 5902 16464 5908 16476
rect 5960 16464 5966 16516
rect 9398 16464 9404 16516
rect 9456 16464 9462 16516
rect 9674 16464 9680 16516
rect 9732 16504 9738 16516
rect 11698 16504 11704 16516
rect 9732 16476 9890 16504
rect 10704 16476 11704 16504
rect 9732 16464 9738 16476
rect 4617 16439 4675 16445
rect 4617 16436 4629 16439
rect 4080 16408 4629 16436
rect 4617 16405 4629 16408
rect 4663 16405 4675 16439
rect 4617 16399 4675 16405
rect 8202 16396 8208 16448
rect 8260 16436 8266 16448
rect 10704 16436 10732 16476
rect 11698 16464 11704 16476
rect 11756 16464 11762 16516
rect 15856 16504 15884 16532
rect 16761 16507 16819 16513
rect 16761 16504 16773 16507
rect 15686 16476 15792 16504
rect 15856 16476 16773 16504
rect 8260 16408 10732 16436
rect 10873 16439 10931 16445
rect 8260 16396 8266 16408
rect 10873 16405 10885 16439
rect 10919 16436 10931 16439
rect 11054 16436 11060 16448
rect 10919 16408 11060 16436
rect 10919 16405 10931 16408
rect 10873 16399 10931 16405
rect 11054 16396 11060 16408
rect 11112 16436 11118 16448
rect 12250 16436 12256 16448
rect 11112 16408 12256 16436
rect 11112 16396 11118 16408
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 15562 16436 15568 16448
rect 13872 16408 15568 16436
rect 13872 16396 13878 16408
rect 15562 16396 15568 16408
rect 15620 16396 15626 16448
rect 15764 16436 15792 16476
rect 16761 16473 16773 16476
rect 16807 16473 16819 16507
rect 17880 16504 17908 16612
rect 17954 16532 17960 16584
rect 18012 16532 18018 16584
rect 18248 16581 18276 16748
rect 19334 16736 19340 16748
rect 19392 16736 19398 16788
rect 20990 16776 20996 16788
rect 20272 16748 20996 16776
rect 18414 16640 18420 16652
rect 18340 16612 18420 16640
rect 18340 16581 18368 16612
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 18233 16575 18291 16581
rect 18233 16541 18245 16575
rect 18279 16541 18291 16575
rect 18233 16535 18291 16541
rect 18325 16575 18383 16581
rect 18325 16541 18337 16575
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 18598 16532 18604 16584
rect 18656 16532 18662 16584
rect 20272 16581 20300 16748
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 29178 16736 29184 16788
rect 29236 16776 29242 16788
rect 30101 16779 30159 16785
rect 30101 16776 30113 16779
rect 29236 16748 30113 16776
rect 29236 16736 29242 16748
rect 30101 16745 30113 16748
rect 30147 16745 30159 16779
rect 30101 16739 30159 16745
rect 31202 16736 31208 16788
rect 31260 16736 31266 16788
rect 32122 16736 32128 16788
rect 32180 16776 32186 16788
rect 32582 16776 32588 16788
rect 32180 16748 32588 16776
rect 32180 16736 32186 16748
rect 32582 16736 32588 16748
rect 32640 16736 32646 16788
rect 35161 16779 35219 16785
rect 35161 16745 35173 16779
rect 35207 16776 35219 16779
rect 35250 16776 35256 16788
rect 35207 16748 35256 16776
rect 35207 16745 35219 16748
rect 35161 16739 35219 16745
rect 35250 16736 35256 16748
rect 35308 16736 35314 16788
rect 35434 16736 35440 16788
rect 35492 16736 35498 16788
rect 20438 16668 20444 16720
rect 20496 16668 20502 16720
rect 20714 16668 20720 16720
rect 20772 16668 20778 16720
rect 25406 16708 25412 16720
rect 23508 16680 25412 16708
rect 20456 16640 20484 16668
rect 20732 16640 20760 16668
rect 20456 16612 20668 16640
rect 20732 16612 21404 16640
rect 20257 16575 20315 16581
rect 20257 16572 20269 16575
rect 18708 16544 20269 16572
rect 18708 16504 18736 16544
rect 20257 16541 20269 16544
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 20346 16532 20352 16584
rect 20404 16572 20410 16584
rect 20640 16581 20668 16612
rect 20806 16581 20812 16584
rect 20625 16575 20683 16581
rect 20404 16544 20449 16572
rect 20404 16532 20410 16544
rect 20625 16541 20637 16575
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 20763 16575 20812 16581
rect 20763 16541 20775 16575
rect 20809 16541 20812 16575
rect 20763 16535 20812 16541
rect 20806 16532 20812 16535
rect 20864 16532 20870 16584
rect 20990 16532 20996 16584
rect 21048 16532 21054 16584
rect 21376 16581 21404 16612
rect 23198 16600 23204 16652
rect 23256 16600 23262 16652
rect 23508 16649 23536 16680
rect 25406 16668 25412 16680
rect 25464 16668 25470 16720
rect 29362 16668 29368 16720
rect 29420 16708 29426 16720
rect 34333 16711 34391 16717
rect 34333 16708 34345 16711
rect 29420 16680 34345 16708
rect 29420 16668 29426 16680
rect 34333 16677 34345 16680
rect 34379 16677 34391 16711
rect 34333 16671 34391 16677
rect 34425 16711 34483 16717
rect 34425 16677 34437 16711
rect 34471 16708 34483 16711
rect 35345 16711 35403 16717
rect 35345 16708 35357 16711
rect 34471 16680 35357 16708
rect 34471 16677 34483 16680
rect 34425 16671 34483 16677
rect 35345 16677 35357 16680
rect 35391 16708 35403 16711
rect 35391 16680 35664 16708
rect 35391 16677 35403 16680
rect 35345 16671 35403 16677
rect 23493 16643 23551 16649
rect 23493 16640 23505 16643
rect 23308 16612 23505 16640
rect 21361 16575 21419 16581
rect 21361 16541 21373 16575
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 21821 16575 21879 16581
rect 21821 16541 21833 16575
rect 21867 16541 21879 16575
rect 21821 16535 21879 16541
rect 17880 16476 18736 16504
rect 16761 16467 16819 16473
rect 19058 16464 19064 16516
rect 19116 16464 19122 16516
rect 20533 16507 20591 16513
rect 20533 16473 20545 16507
rect 20579 16473 20591 16507
rect 21836 16504 21864 16535
rect 22278 16532 22284 16584
rect 22336 16532 22342 16584
rect 22922 16572 22928 16584
rect 22388 16544 22928 16572
rect 22388 16516 22416 16544
rect 22922 16532 22928 16544
rect 22980 16532 22986 16584
rect 23308 16572 23336 16612
rect 23493 16609 23505 16612
rect 23539 16609 23551 16643
rect 23493 16603 23551 16609
rect 23937 16643 23995 16649
rect 23937 16609 23949 16643
rect 23983 16640 23995 16643
rect 24854 16640 24860 16652
rect 23983 16612 24860 16640
rect 23983 16609 23995 16612
rect 23937 16603 23995 16609
rect 24854 16600 24860 16612
rect 24912 16640 24918 16652
rect 25593 16643 25651 16649
rect 24912 16612 25544 16640
rect 24912 16600 24918 16612
rect 23216 16544 23336 16572
rect 23216 16516 23244 16544
rect 23382 16532 23388 16584
rect 23440 16532 23446 16584
rect 25222 16532 25228 16584
rect 25280 16532 25286 16584
rect 25409 16575 25467 16581
rect 25409 16541 25421 16575
rect 25455 16541 25467 16575
rect 25516 16572 25544 16612
rect 25593 16609 25605 16643
rect 25639 16640 25651 16643
rect 26234 16640 26240 16652
rect 25639 16612 26240 16640
rect 25639 16609 25651 16612
rect 25593 16603 25651 16609
rect 26234 16600 26240 16612
rect 26292 16600 26298 16652
rect 32582 16640 32588 16652
rect 30024 16612 32588 16640
rect 26050 16572 26056 16584
rect 25516 16544 26056 16572
rect 25409 16535 25467 16541
rect 20533 16467 20591 16473
rect 20916 16476 21864 16504
rect 22097 16507 22155 16513
rect 16298 16436 16304 16448
rect 15764 16408 16304 16436
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 16390 16396 16396 16448
rect 16448 16436 16454 16448
rect 16485 16439 16543 16445
rect 16485 16436 16497 16439
rect 16448 16408 16497 16436
rect 16448 16396 16454 16408
rect 16485 16405 16497 16408
rect 16531 16405 16543 16439
rect 16485 16399 16543 16405
rect 16942 16396 16948 16448
rect 17000 16436 17006 16448
rect 17129 16439 17187 16445
rect 17129 16436 17141 16439
rect 17000 16408 17141 16436
rect 17000 16396 17006 16408
rect 17129 16405 17141 16408
rect 17175 16405 17187 16439
rect 17129 16399 17187 16405
rect 18138 16396 18144 16448
rect 18196 16436 18202 16448
rect 18506 16436 18512 16448
rect 18196 16408 18512 16436
rect 18196 16396 18202 16408
rect 18506 16396 18512 16408
rect 18564 16436 18570 16448
rect 20548 16436 20576 16467
rect 20916 16448 20944 16476
rect 22097 16473 22109 16507
rect 22143 16504 22155 16507
rect 22370 16504 22376 16516
rect 22143 16476 22376 16504
rect 22143 16473 22155 16476
rect 22097 16467 22155 16473
rect 22370 16464 22376 16476
rect 22428 16464 22434 16516
rect 22830 16464 22836 16516
rect 22888 16464 22894 16516
rect 23198 16464 23204 16516
rect 23256 16464 23262 16516
rect 23290 16464 23296 16516
rect 23348 16464 23354 16516
rect 18564 16408 20576 16436
rect 18564 16396 18570 16408
rect 20898 16396 20904 16448
rect 20956 16396 20962 16448
rect 23400 16445 23428 16532
rect 23750 16464 23756 16516
rect 23808 16464 23814 16516
rect 25424 16504 25452 16535
rect 26050 16532 26056 16544
rect 26108 16532 26114 16584
rect 30024 16581 30052 16612
rect 32582 16600 32588 16612
rect 32640 16600 32646 16652
rect 34241 16643 34299 16649
rect 34241 16609 34253 16643
rect 34287 16640 34299 16643
rect 35526 16640 35532 16652
rect 34287 16612 35532 16640
rect 34287 16609 34299 16612
rect 34241 16603 34299 16609
rect 35526 16600 35532 16612
rect 35584 16600 35590 16652
rect 30009 16575 30067 16581
rect 30009 16541 30021 16575
rect 30055 16541 30067 16575
rect 30009 16535 30067 16541
rect 30190 16532 30196 16584
rect 30248 16532 30254 16584
rect 30282 16532 30288 16584
rect 30340 16572 30346 16584
rect 30561 16575 30619 16581
rect 30561 16572 30573 16575
rect 30340 16544 30573 16572
rect 30340 16532 30346 16544
rect 30561 16541 30573 16544
rect 30607 16541 30619 16575
rect 30561 16535 30619 16541
rect 30650 16532 30656 16584
rect 30708 16572 30714 16584
rect 30745 16575 30803 16581
rect 30745 16572 30757 16575
rect 30708 16544 30757 16572
rect 30708 16532 30714 16544
rect 30745 16541 30757 16544
rect 30791 16572 30803 16575
rect 30926 16572 30932 16584
rect 30791 16544 30932 16572
rect 30791 16541 30803 16544
rect 30745 16535 30803 16541
rect 30926 16532 30932 16544
rect 30984 16532 30990 16584
rect 31389 16575 31447 16581
rect 31389 16541 31401 16575
rect 31435 16572 31447 16575
rect 31478 16572 31484 16584
rect 31435 16544 31484 16572
rect 31435 16541 31447 16544
rect 31389 16535 31447 16541
rect 31478 16532 31484 16544
rect 31536 16532 31542 16584
rect 31754 16532 31760 16584
rect 31812 16572 31818 16584
rect 32309 16575 32367 16581
rect 32309 16572 32321 16575
rect 31812 16544 32321 16572
rect 31812 16532 31818 16544
rect 32309 16541 32321 16544
rect 32355 16541 32367 16575
rect 35437 16575 35495 16581
rect 32309 16535 32367 16541
rect 34516 16553 34574 16559
rect 34516 16519 34528 16553
rect 34562 16519 34574 16553
rect 35437 16541 35449 16575
rect 35483 16572 35495 16575
rect 35636 16572 35664 16680
rect 35483 16544 35664 16572
rect 35483 16541 35495 16544
rect 35437 16535 35495 16541
rect 34516 16516 34574 16519
rect 25148 16476 25452 16504
rect 25148 16448 25176 16476
rect 25498 16464 25504 16516
rect 25556 16504 25562 16516
rect 26237 16507 26295 16513
rect 26237 16504 26249 16507
rect 25556 16476 26249 16504
rect 25556 16464 25562 16476
rect 26237 16473 26249 16476
rect 26283 16473 26295 16507
rect 26237 16467 26295 16473
rect 29270 16464 29276 16516
rect 29328 16504 29334 16516
rect 29328 16476 31754 16504
rect 29328 16464 29334 16476
rect 23385 16439 23443 16445
rect 23385 16405 23397 16439
rect 23431 16405 23443 16439
rect 23385 16399 23443 16405
rect 25130 16396 25136 16448
rect 25188 16396 25194 16448
rect 26418 16396 26424 16448
rect 26476 16396 26482 16448
rect 28074 16396 28080 16448
rect 28132 16436 28138 16448
rect 30650 16436 30656 16448
rect 28132 16408 30656 16436
rect 28132 16396 28138 16408
rect 30650 16396 30656 16408
rect 30708 16396 30714 16448
rect 30742 16396 30748 16448
rect 30800 16396 30806 16448
rect 31726 16436 31754 16476
rect 32490 16464 32496 16516
rect 32548 16464 32554 16516
rect 34514 16464 34520 16516
rect 34572 16464 34578 16516
rect 34790 16464 34796 16516
rect 34848 16504 34854 16516
rect 34977 16507 35035 16513
rect 34977 16504 34989 16507
rect 34848 16476 34989 16504
rect 34848 16464 34854 16476
rect 34977 16473 34989 16476
rect 35023 16473 35035 16507
rect 34977 16467 35035 16473
rect 35084 16476 35848 16504
rect 35084 16436 35112 16476
rect 31726 16408 35112 16436
rect 35158 16396 35164 16448
rect 35216 16445 35222 16448
rect 35820 16445 35848 16476
rect 35216 16439 35235 16445
rect 35223 16405 35235 16439
rect 35216 16399 35235 16405
rect 35805 16439 35863 16445
rect 35805 16405 35817 16439
rect 35851 16405 35863 16439
rect 35805 16399 35863 16405
rect 35216 16396 35222 16399
rect 1104 16346 38272 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38272 16346
rect 1104 16272 38272 16294
rect 1394 16192 1400 16244
rect 1452 16232 1458 16244
rect 2958 16232 2964 16244
rect 1452 16204 2964 16232
rect 1452 16192 1458 16204
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 3602 16192 3608 16244
rect 3660 16232 3666 16244
rect 3881 16235 3939 16241
rect 3881 16232 3893 16235
rect 3660 16204 3893 16232
rect 3660 16192 3666 16204
rect 3881 16201 3893 16204
rect 3927 16201 3939 16235
rect 3881 16195 3939 16201
rect 4049 16235 4107 16241
rect 4049 16201 4061 16235
rect 4095 16232 4107 16235
rect 4614 16232 4620 16244
rect 4095 16204 4620 16232
rect 4095 16201 4107 16204
rect 4049 16195 4107 16201
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5169 16235 5227 16241
rect 5169 16232 5181 16235
rect 5040 16204 5181 16232
rect 5040 16192 5046 16204
rect 5169 16201 5181 16204
rect 5215 16201 5227 16235
rect 5442 16232 5448 16244
rect 5169 16195 5227 16201
rect 5368 16204 5448 16232
rect 1673 16167 1731 16173
rect 1673 16133 1685 16167
rect 1719 16164 1731 16167
rect 1946 16164 1952 16176
rect 1719 16136 1952 16164
rect 1719 16133 1731 16136
rect 1673 16127 1731 16133
rect 1946 16124 1952 16136
rect 2004 16124 2010 16176
rect 4249 16167 4307 16173
rect 4249 16133 4261 16167
rect 4295 16164 4307 16167
rect 4798 16164 4804 16176
rect 4295 16136 4804 16164
rect 4295 16133 4307 16136
rect 4249 16127 4307 16133
rect 4798 16124 4804 16136
rect 4856 16124 4862 16176
rect 5368 16096 5396 16204
rect 5442 16192 5448 16204
rect 5500 16192 5506 16244
rect 9398 16192 9404 16244
rect 9456 16232 9462 16244
rect 9493 16235 9551 16241
rect 9493 16232 9505 16235
rect 9456 16204 9505 16232
rect 9456 16192 9462 16204
rect 9493 16201 9505 16204
rect 9539 16201 9551 16235
rect 9493 16195 9551 16201
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16201 9827 16235
rect 9769 16195 9827 16201
rect 10137 16235 10195 16241
rect 10137 16201 10149 16235
rect 10183 16232 10195 16235
rect 12526 16232 12532 16244
rect 10183 16204 12532 16232
rect 10183 16201 10195 16204
rect 10137 16195 10195 16201
rect 2806 16068 5396 16096
rect 5460 16136 6040 16164
rect 1394 15988 1400 16040
rect 1452 15988 1458 16040
rect 2130 15988 2136 16040
rect 2188 16028 2194 16040
rect 5460 16028 5488 16136
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16065 5595 16099
rect 5537 16059 5595 16065
rect 2188 16000 5488 16028
rect 2188 15988 2194 16000
rect 5552 15960 5580 16059
rect 5626 15988 5632 16040
rect 5684 15988 5690 16040
rect 5813 16031 5871 16037
rect 5813 15997 5825 16031
rect 5859 16028 5871 16031
rect 5902 16028 5908 16040
rect 5859 16000 5908 16028
rect 5859 15997 5871 16000
rect 5813 15991 5871 15997
rect 5902 15988 5908 16000
rect 5960 15988 5966 16040
rect 6012 16028 6040 16136
rect 9677 16099 9735 16105
rect 9677 16065 9689 16099
rect 9723 16096 9735 16099
rect 9784 16096 9812 16195
rect 12526 16192 12532 16204
rect 12584 16232 12590 16244
rect 13170 16232 13176 16244
rect 12584 16204 13176 16232
rect 12584 16192 12590 16204
rect 13170 16192 13176 16204
rect 13228 16192 13234 16244
rect 14458 16192 14464 16244
rect 14516 16192 14522 16244
rect 14550 16192 14556 16244
rect 14608 16232 14614 16244
rect 16390 16232 16396 16244
rect 14608 16204 16396 16232
rect 14608 16192 14614 16204
rect 16390 16192 16396 16204
rect 16448 16192 16454 16244
rect 16850 16192 16856 16244
rect 16908 16192 16914 16244
rect 17310 16192 17316 16244
rect 17368 16232 17374 16244
rect 17697 16235 17755 16241
rect 17697 16232 17709 16235
rect 17368 16204 17709 16232
rect 17368 16192 17374 16204
rect 17697 16201 17709 16204
rect 17743 16201 17755 16235
rect 17697 16195 17755 16201
rect 17865 16235 17923 16241
rect 17865 16201 17877 16235
rect 17911 16201 17923 16235
rect 17865 16195 17923 16201
rect 10229 16167 10287 16173
rect 10229 16133 10241 16167
rect 10275 16164 10287 16167
rect 11054 16164 11060 16176
rect 10275 16136 11060 16164
rect 10275 16133 10287 16136
rect 10229 16127 10287 16133
rect 11054 16124 11060 16136
rect 11112 16124 11118 16176
rect 12986 16124 12992 16176
rect 13044 16164 13050 16176
rect 17218 16164 17224 16176
rect 13044 16136 17224 16164
rect 13044 16124 13050 16136
rect 17218 16124 17224 16136
rect 17276 16164 17282 16176
rect 17497 16167 17555 16173
rect 17497 16164 17509 16167
rect 17276 16136 17509 16164
rect 17276 16124 17282 16136
rect 17497 16133 17509 16136
rect 17543 16164 17555 16167
rect 17880 16164 17908 16195
rect 19058 16192 19064 16244
rect 19116 16192 19122 16244
rect 19426 16192 19432 16244
rect 19484 16192 19490 16244
rect 20272 16204 20668 16232
rect 18785 16167 18843 16173
rect 18785 16164 18797 16167
rect 17543 16136 17816 16164
rect 17880 16136 18797 16164
rect 17543 16133 17555 16136
rect 17497 16127 17555 16133
rect 9723 16068 9812 16096
rect 9876 16068 11284 16096
rect 9723 16065 9735 16068
rect 9677 16059 9735 16065
rect 9876 16028 9904 16068
rect 11256 16040 11284 16068
rect 12250 16056 12256 16108
rect 12308 16056 12314 16108
rect 12342 16056 12348 16108
rect 12400 16056 12406 16108
rect 14001 16099 14059 16105
rect 14001 16065 14013 16099
rect 14047 16096 14059 16099
rect 14182 16096 14188 16108
rect 14047 16068 14188 16096
rect 14047 16065 14059 16068
rect 14001 16059 14059 16065
rect 14182 16056 14188 16068
rect 14240 16056 14246 16108
rect 14277 16099 14335 16105
rect 14277 16065 14289 16099
rect 14323 16096 14335 16099
rect 14550 16096 14556 16108
rect 14323 16068 14556 16096
rect 14323 16065 14335 16068
rect 14277 16059 14335 16065
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 16390 16056 16396 16108
rect 16448 16096 16454 16108
rect 16945 16099 17003 16105
rect 16945 16096 16957 16099
rect 16448 16068 16957 16096
rect 16448 16056 16454 16068
rect 16945 16065 16957 16068
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 17034 16056 17040 16108
rect 17092 16056 17098 16108
rect 17788 16096 17816 16136
rect 18785 16133 18797 16136
rect 18831 16133 18843 16167
rect 18785 16127 18843 16133
rect 17957 16099 18015 16105
rect 17957 16096 17969 16099
rect 17788 16068 17969 16096
rect 17957 16065 17969 16068
rect 18003 16065 18015 16099
rect 17957 16059 18015 16065
rect 18138 16056 18144 16108
rect 18196 16056 18202 16108
rect 18230 16056 18236 16108
rect 18288 16056 18294 16108
rect 18322 16056 18328 16108
rect 18380 16096 18386 16108
rect 18874 16096 18880 16108
rect 18380 16068 18880 16096
rect 18380 16056 18386 16068
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 6012 16000 9904 16028
rect 10318 15988 10324 16040
rect 10376 15988 10382 16040
rect 11238 15988 11244 16040
rect 11296 15988 11302 16040
rect 11606 15988 11612 16040
rect 11664 16028 11670 16040
rect 12529 16031 12587 16037
rect 12529 16028 12541 16031
rect 11664 16000 12541 16028
rect 11664 15988 11670 16000
rect 12529 15997 12541 16000
rect 12575 16028 12587 16031
rect 17052 16028 17080 16056
rect 12575 16000 16988 16028
rect 17052 16000 19012 16028
rect 12575 15997 12587 16000
rect 12529 15991 12587 15997
rect 11885 15963 11943 15969
rect 11885 15960 11897 15963
rect 5552 15932 11897 15960
rect 11885 15929 11897 15932
rect 11931 15929 11943 15963
rect 11885 15923 11943 15929
rect 12158 15920 12164 15972
rect 12216 15960 12222 15972
rect 13354 15960 13360 15972
rect 12216 15932 13360 15960
rect 12216 15920 12222 15932
rect 13354 15920 13360 15932
rect 13412 15920 13418 15972
rect 14093 15963 14151 15969
rect 14093 15929 14105 15963
rect 14139 15960 14151 15963
rect 15102 15960 15108 15972
rect 14139 15932 15108 15960
rect 14139 15929 14151 15932
rect 14093 15923 14151 15929
rect 15102 15920 15108 15932
rect 15160 15920 15166 15972
rect 16850 15960 16856 15972
rect 16592 15932 16856 15960
rect 3142 15852 3148 15904
rect 3200 15892 3206 15904
rect 3878 15892 3884 15904
rect 3200 15864 3884 15892
rect 3200 15852 3206 15864
rect 3878 15852 3884 15864
rect 3936 15892 3942 15904
rect 4065 15895 4123 15901
rect 4065 15892 4077 15895
rect 3936 15864 4077 15892
rect 3936 15852 3942 15864
rect 4065 15861 4077 15864
rect 4111 15892 4123 15895
rect 16592 15892 16620 15932
rect 16850 15920 16856 15932
rect 16908 15920 16914 15972
rect 4111 15864 16620 15892
rect 4111 15861 4123 15864
rect 4065 15855 4123 15861
rect 16666 15852 16672 15904
rect 16724 15852 16730 15904
rect 16960 15892 16988 16000
rect 17126 15920 17132 15972
rect 17184 15960 17190 15972
rect 17221 15963 17279 15969
rect 17221 15960 17233 15963
rect 17184 15932 17233 15960
rect 17184 15920 17190 15932
rect 17221 15929 17233 15932
rect 17267 15929 17279 15963
rect 17221 15923 17279 15929
rect 17328 15932 18736 15960
rect 17328 15892 17356 15932
rect 18708 15904 18736 15932
rect 16960 15864 17356 15892
rect 17681 15895 17739 15901
rect 17681 15861 17693 15895
rect 17727 15892 17739 15895
rect 18322 15892 18328 15904
rect 17727 15864 18328 15892
rect 17727 15861 17739 15864
rect 17681 15855 17739 15861
rect 18322 15852 18328 15864
rect 18380 15852 18386 15904
rect 18598 15852 18604 15904
rect 18656 15852 18662 15904
rect 18690 15852 18696 15904
rect 18748 15892 18754 15904
rect 18877 15895 18935 15901
rect 18877 15892 18889 15895
rect 18748 15864 18889 15892
rect 18748 15852 18754 15864
rect 18877 15861 18889 15864
rect 18923 15861 18935 15895
rect 18984 15892 19012 16000
rect 19076 15960 19104 16192
rect 19444 16096 19472 16192
rect 20272 16105 20300 16204
rect 20349 16167 20407 16173
rect 20349 16133 20361 16167
rect 20395 16164 20407 16167
rect 20438 16164 20444 16176
rect 20395 16136 20444 16164
rect 20395 16133 20407 16136
rect 20349 16127 20407 16133
rect 20438 16124 20444 16136
rect 20496 16124 20502 16176
rect 20549 16167 20607 16173
rect 20549 16133 20561 16167
rect 20595 16133 20607 16167
rect 20549 16127 20607 16133
rect 20257 16099 20315 16105
rect 20257 16096 20269 16099
rect 19444 16068 20269 16096
rect 20257 16065 20269 16068
rect 20303 16065 20315 16099
rect 20257 16059 20315 16065
rect 20564 16040 20592 16127
rect 20640 16040 20668 16204
rect 20714 16192 20720 16244
rect 20772 16192 20778 16244
rect 20806 16192 20812 16244
rect 20864 16232 20870 16244
rect 21266 16232 21272 16244
rect 20864 16204 21272 16232
rect 20864 16192 20870 16204
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 21453 16235 21511 16241
rect 21453 16201 21465 16235
rect 21499 16232 21511 16235
rect 22278 16232 22284 16244
rect 21499 16204 22284 16232
rect 21499 16201 21511 16204
rect 21453 16195 21511 16201
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 25222 16192 25228 16244
rect 25280 16232 25286 16244
rect 25280 16204 26372 16232
rect 25280 16192 25286 16204
rect 23014 16124 23020 16176
rect 23072 16124 23078 16176
rect 25130 16124 25136 16176
rect 25188 16164 25194 16176
rect 25188 16136 26280 16164
rect 25188 16124 25194 16136
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21269 16099 21327 16105
rect 21269 16096 21281 16099
rect 20956 16068 21281 16096
rect 20956 16056 20962 16068
rect 21269 16065 21281 16068
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 21450 16056 21456 16108
rect 21508 16096 21514 16108
rect 22002 16096 22008 16108
rect 21508 16068 22008 16096
rect 21508 16056 21514 16068
rect 22002 16056 22008 16068
rect 22060 16096 22066 16108
rect 22833 16099 22891 16105
rect 22833 16096 22845 16099
rect 22060 16068 22845 16096
rect 22060 16056 22066 16068
rect 22833 16065 22845 16068
rect 22879 16065 22891 16099
rect 22833 16059 22891 16065
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16065 23167 16099
rect 23109 16059 23167 16065
rect 20530 15988 20536 16040
rect 20588 15988 20594 16040
rect 20622 15988 20628 16040
rect 20680 15988 20686 16040
rect 20806 15988 20812 16040
rect 20864 16028 20870 16040
rect 20990 16028 20996 16040
rect 20864 16000 20996 16028
rect 20864 15988 20870 16000
rect 20990 15988 20996 16000
rect 21048 15988 21054 16040
rect 21358 15988 21364 16040
rect 21416 16028 21422 16040
rect 23124 16028 23152 16059
rect 23198 16056 23204 16108
rect 23256 16056 23262 16108
rect 24670 16056 24676 16108
rect 24728 16056 24734 16108
rect 24854 16056 24860 16108
rect 24912 16096 24918 16108
rect 26252 16105 26280 16136
rect 26344 16105 26372 16204
rect 29178 16192 29184 16244
rect 29236 16232 29242 16244
rect 29273 16235 29331 16241
rect 29273 16232 29285 16235
rect 29236 16204 29285 16232
rect 29236 16192 29242 16204
rect 29273 16201 29285 16204
rect 29319 16201 29331 16235
rect 29273 16195 29331 16201
rect 30190 16192 30196 16244
rect 30248 16232 30254 16244
rect 30469 16235 30527 16241
rect 30469 16232 30481 16235
rect 30248 16204 30481 16232
rect 30248 16192 30254 16204
rect 30469 16201 30481 16204
rect 30515 16201 30527 16235
rect 30469 16195 30527 16201
rect 30742 16192 30748 16244
rect 30800 16232 30806 16244
rect 30837 16235 30895 16241
rect 30837 16232 30849 16235
rect 30800 16204 30849 16232
rect 30800 16192 30806 16204
rect 30837 16201 30849 16204
rect 30883 16201 30895 16235
rect 30837 16195 30895 16201
rect 30926 16192 30932 16244
rect 30984 16232 30990 16244
rect 30984 16204 31248 16232
rect 30984 16192 30990 16204
rect 29383 16167 29441 16173
rect 29383 16164 29395 16167
rect 27264 16136 27614 16164
rect 25225 16099 25283 16105
rect 25225 16096 25237 16099
rect 24912 16068 25237 16096
rect 24912 16056 24918 16068
rect 25225 16065 25237 16068
rect 25271 16065 25283 16099
rect 25225 16059 25283 16065
rect 26237 16099 26295 16105
rect 26237 16065 26249 16099
rect 26283 16065 26295 16099
rect 26237 16059 26295 16065
rect 26329 16099 26387 16105
rect 26329 16065 26341 16099
rect 26375 16065 26387 16099
rect 26329 16059 26387 16065
rect 26418 16056 26424 16108
rect 26476 16096 26482 16108
rect 27065 16099 27123 16105
rect 27065 16096 27077 16099
rect 26476 16068 27077 16096
rect 26476 16056 26482 16068
rect 27065 16065 27077 16068
rect 27111 16065 27123 16099
rect 27065 16059 27123 16065
rect 27264 16037 27292 16136
rect 27341 16099 27399 16105
rect 27341 16065 27353 16099
rect 27387 16065 27399 16099
rect 27341 16059 27399 16065
rect 21416 16000 23152 16028
rect 26513 16031 26571 16037
rect 21416 15988 21422 16000
rect 26513 15997 26525 16031
rect 26559 16028 26571 16031
rect 27249 16031 27307 16037
rect 27249 16028 27261 16031
rect 26559 16000 27261 16028
rect 26559 15997 26571 16000
rect 26513 15991 26571 15997
rect 27249 15997 27261 16000
rect 27295 15997 27307 16031
rect 27249 15991 27307 15997
rect 27356 15972 27384 16059
rect 27586 16028 27614 16136
rect 29104 16136 29395 16164
rect 29104 16108 29132 16136
rect 29383 16133 29395 16136
rect 29429 16133 29441 16167
rect 29549 16167 29607 16173
rect 29549 16164 29561 16167
rect 29383 16127 29441 16133
rect 29472 16136 29561 16164
rect 29086 16056 29092 16108
rect 29144 16056 29150 16108
rect 29264 16099 29322 16105
rect 29264 16096 29276 16099
rect 29196 16068 29276 16096
rect 29196 16028 29224 16068
rect 29264 16065 29276 16068
rect 29310 16065 29322 16099
rect 29264 16059 29322 16065
rect 29472 16040 29500 16136
rect 29549 16133 29561 16136
rect 29595 16133 29607 16167
rect 29549 16127 29607 16133
rect 29638 16124 29644 16176
rect 29696 16164 29702 16176
rect 30282 16164 30288 16176
rect 29696 16136 30288 16164
rect 29696 16124 29702 16136
rect 30116 16105 30144 16136
rect 30282 16124 30288 16136
rect 30340 16164 30346 16176
rect 31220 16173 31248 16204
rect 34790 16192 34796 16244
rect 34848 16232 34854 16244
rect 34977 16235 35035 16241
rect 34977 16232 34989 16235
rect 34848 16204 34989 16232
rect 34848 16192 34854 16204
rect 34977 16201 34989 16204
rect 35023 16201 35035 16235
rect 34977 16195 35035 16201
rect 35250 16192 35256 16244
rect 35308 16192 35314 16244
rect 31021 16167 31079 16173
rect 31021 16164 31033 16167
rect 30340 16136 31033 16164
rect 30340 16124 30346 16136
rect 31021 16133 31033 16136
rect 31067 16133 31079 16167
rect 31021 16127 31079 16133
rect 31205 16167 31263 16173
rect 31205 16133 31217 16167
rect 31251 16133 31263 16167
rect 35268 16164 35296 16192
rect 31205 16127 31263 16133
rect 34900 16136 35296 16164
rect 34900 16105 34928 16136
rect 30101 16099 30159 16105
rect 30101 16065 30113 16099
rect 30147 16065 30159 16099
rect 30101 16059 30159 16065
rect 30653 16099 30711 16105
rect 30653 16065 30665 16099
rect 30699 16065 30711 16099
rect 30653 16059 30711 16065
rect 30929 16099 30987 16105
rect 30929 16065 30941 16099
rect 30975 16065 30987 16099
rect 30929 16059 30987 16065
rect 34885 16099 34943 16105
rect 34885 16065 34897 16099
rect 34931 16065 34943 16099
rect 34885 16059 34943 16065
rect 29454 16028 29460 16040
rect 27586 16000 29460 16028
rect 29454 15988 29460 16000
rect 29512 15988 29518 16040
rect 29733 16031 29791 16037
rect 29733 15997 29745 16031
rect 29779 16028 29791 16031
rect 29917 16031 29975 16037
rect 29917 16028 29929 16031
rect 29779 16000 29929 16028
rect 29779 15997 29791 16000
rect 29733 15991 29791 15997
rect 29917 15997 29929 16000
rect 29963 15997 29975 16031
rect 29917 15991 29975 15997
rect 27154 15960 27160 15972
rect 19076 15932 27160 15960
rect 27154 15920 27160 15932
rect 27212 15920 27218 15972
rect 27338 15920 27344 15972
rect 27396 15960 27402 15972
rect 30668 15960 30696 16059
rect 30944 16028 30972 16059
rect 35158 16056 35164 16108
rect 35216 16056 35222 16108
rect 37645 16099 37703 16105
rect 37645 16065 37657 16099
rect 37691 16065 37703 16099
rect 37645 16059 37703 16065
rect 32214 16028 32220 16040
rect 30944 16000 32220 16028
rect 32214 15988 32220 16000
rect 32272 15988 32278 16040
rect 34790 15988 34796 16040
rect 34848 16028 34854 16040
rect 35176 16028 35204 16056
rect 34848 16000 35204 16028
rect 34848 15988 34854 16000
rect 37660 15960 37688 16059
rect 27396 15932 30696 15960
rect 30760 15932 37688 15960
rect 27396 15920 27402 15932
rect 20165 15895 20223 15901
rect 20165 15892 20177 15895
rect 18984 15864 20177 15892
rect 18877 15855 18935 15861
rect 20165 15861 20177 15864
rect 20211 15861 20223 15895
rect 20165 15855 20223 15861
rect 20438 15852 20444 15904
rect 20496 15892 20502 15904
rect 20533 15895 20591 15901
rect 20533 15892 20545 15895
rect 20496 15864 20545 15892
rect 20496 15852 20502 15864
rect 20533 15861 20545 15864
rect 20579 15861 20591 15895
rect 20533 15855 20591 15861
rect 20714 15852 20720 15904
rect 20772 15892 20778 15904
rect 21085 15895 21143 15901
rect 21085 15892 21097 15895
rect 20772 15864 21097 15892
rect 20772 15852 20778 15864
rect 21085 15861 21097 15864
rect 21131 15861 21143 15895
rect 21085 15855 21143 15861
rect 23385 15895 23443 15901
rect 23385 15861 23397 15895
rect 23431 15892 23443 15895
rect 24946 15892 24952 15904
rect 23431 15864 24952 15892
rect 23431 15861 23443 15864
rect 23385 15855 23443 15861
rect 24946 15852 24952 15864
rect 25004 15852 25010 15904
rect 25038 15852 25044 15904
rect 25096 15892 25102 15904
rect 25685 15895 25743 15901
rect 25685 15892 25697 15895
rect 25096 15864 25697 15892
rect 25096 15852 25102 15864
rect 25685 15861 25697 15864
rect 25731 15892 25743 15895
rect 27430 15892 27436 15904
rect 25731 15864 27436 15892
rect 25731 15861 25743 15864
rect 25685 15855 25743 15861
rect 27430 15852 27436 15864
rect 27488 15852 27494 15904
rect 27525 15895 27583 15901
rect 27525 15861 27537 15895
rect 27571 15892 27583 15895
rect 29362 15892 29368 15904
rect 27571 15864 29368 15892
rect 27571 15861 27583 15864
rect 27525 15855 27583 15861
rect 29362 15852 29368 15864
rect 29420 15852 29426 15904
rect 30098 15852 30104 15904
rect 30156 15892 30162 15904
rect 30285 15895 30343 15901
rect 30285 15892 30297 15895
rect 30156 15864 30297 15892
rect 30156 15852 30162 15864
rect 30285 15861 30297 15864
rect 30331 15861 30343 15895
rect 30285 15855 30343 15861
rect 30374 15852 30380 15904
rect 30432 15892 30438 15904
rect 30760 15892 30788 15932
rect 30432 15864 30788 15892
rect 30432 15852 30438 15864
rect 31386 15852 31392 15904
rect 31444 15852 31450 15904
rect 34514 15852 34520 15904
rect 34572 15892 34578 15904
rect 35161 15895 35219 15901
rect 35161 15892 35173 15895
rect 34572 15864 35173 15892
rect 34572 15852 34578 15864
rect 35161 15861 35173 15864
rect 35207 15892 35219 15895
rect 35250 15892 35256 15904
rect 35207 15864 35256 15892
rect 35207 15861 35219 15864
rect 35161 15855 35219 15861
rect 35250 15852 35256 15864
rect 35308 15852 35314 15904
rect 37826 15852 37832 15904
rect 37884 15852 37890 15904
rect 1104 15802 38272 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38272 15802
rect 1104 15728 38272 15750
rect 934 15648 940 15700
rect 992 15688 998 15700
rect 1489 15691 1547 15697
rect 1489 15688 1501 15691
rect 992 15660 1501 15688
rect 992 15648 998 15660
rect 1489 15657 1501 15660
rect 1535 15657 1547 15691
rect 1489 15651 1547 15657
rect 3789 15691 3847 15697
rect 3789 15657 3801 15691
rect 3835 15688 3847 15691
rect 3970 15688 3976 15700
rect 3835 15660 3976 15688
rect 3835 15657 3847 15660
rect 3789 15651 3847 15657
rect 3970 15648 3976 15660
rect 4028 15648 4034 15700
rect 4706 15648 4712 15700
rect 4764 15648 4770 15700
rect 4985 15691 5043 15697
rect 4985 15657 4997 15691
rect 5031 15688 5043 15691
rect 5626 15688 5632 15700
rect 5031 15660 5632 15688
rect 5031 15657 5043 15660
rect 4985 15651 5043 15657
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 7558 15688 7564 15700
rect 6288 15660 7564 15688
rect 4614 15620 4620 15632
rect 4540 15592 4620 15620
rect 4540 15561 4568 15592
rect 4614 15580 4620 15592
rect 4672 15580 4678 15632
rect 4724 15620 4752 15648
rect 6288 15620 6316 15660
rect 7558 15648 7564 15660
rect 7616 15688 7622 15700
rect 7929 15691 7987 15697
rect 7929 15688 7941 15691
rect 7616 15660 7941 15688
rect 7616 15648 7622 15660
rect 7929 15657 7941 15660
rect 7975 15657 7987 15691
rect 7929 15651 7987 15657
rect 10226 15648 10232 15700
rect 10284 15688 10290 15700
rect 11054 15688 11060 15700
rect 10284 15660 11060 15688
rect 10284 15648 10290 15660
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 14240 15660 14289 15688
rect 14240 15648 14246 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 14918 15688 14924 15700
rect 14783 15660 14924 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 15562 15648 15568 15700
rect 15620 15688 15626 15700
rect 15838 15688 15844 15700
rect 15620 15660 15844 15688
rect 15620 15648 15626 15660
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 16758 15648 16764 15700
rect 16816 15688 16822 15700
rect 18141 15691 18199 15697
rect 18141 15688 18153 15691
rect 16816 15660 18153 15688
rect 16816 15648 16822 15660
rect 18141 15657 18153 15660
rect 18187 15657 18199 15691
rect 23198 15688 23204 15700
rect 18141 15651 18199 15657
rect 18892 15660 23204 15688
rect 11606 15620 11612 15632
rect 4724 15592 6316 15620
rect 11532 15592 11612 15620
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4525 15555 4583 15561
rect 4111 15524 4476 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 1762 15444 1768 15496
rect 1820 15444 1826 15496
rect 3878 15444 3884 15496
rect 3936 15444 3942 15496
rect 3970 15444 3976 15496
rect 4028 15444 4034 15496
rect 4154 15444 4160 15496
rect 4212 15444 4218 15496
rect 4249 15487 4307 15493
rect 4249 15453 4261 15487
rect 4295 15453 4307 15487
rect 4448 15484 4476 15524
rect 4525 15521 4537 15555
rect 4571 15521 4583 15555
rect 4525 15515 4583 15521
rect 6178 15512 6184 15564
rect 6236 15512 6242 15564
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 11532 15561 11560 15592
rect 11606 15580 11612 15592
rect 11664 15580 11670 15632
rect 11517 15555 11575 15561
rect 11517 15552 11529 15555
rect 11296 15524 11529 15552
rect 11296 15512 11302 15524
rect 11517 15521 11529 15524
rect 11563 15521 11575 15555
rect 15473 15555 15531 15561
rect 15473 15552 15485 15555
rect 11517 15515 11575 15521
rect 14200 15524 15485 15552
rect 4617 15487 4675 15493
rect 4617 15484 4629 15487
rect 4448 15456 4629 15484
rect 4249 15447 4307 15453
rect 4617 15453 4629 15456
rect 4663 15484 4675 15487
rect 4798 15484 4804 15496
rect 4663 15456 4804 15484
rect 4663 15453 4675 15456
rect 4617 15447 4675 15453
rect 3896 15416 3924 15444
rect 4264 15416 4292 15447
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 3896 15388 4292 15416
rect 6196 15416 6224 15512
rect 7834 15444 7840 15496
rect 7892 15484 7898 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 7892 15456 8953 15484
rect 7892 15444 7898 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 11330 15444 11336 15496
rect 11388 15444 11394 15496
rect 11882 15444 11888 15496
rect 11940 15444 11946 15496
rect 14200 15493 14228 15524
rect 15473 15521 15485 15524
rect 15519 15521 15531 15555
rect 15473 15515 15531 15521
rect 15746 15512 15752 15564
rect 15804 15512 15810 15564
rect 15856 15561 15884 15648
rect 18892 15632 18920 15660
rect 23198 15648 23204 15660
rect 23256 15648 23262 15700
rect 24486 15648 24492 15700
rect 24544 15688 24550 15700
rect 26329 15691 26387 15697
rect 24544 15660 25452 15688
rect 24544 15648 24550 15660
rect 17678 15620 17684 15632
rect 16040 15592 17684 15620
rect 15841 15555 15899 15561
rect 15841 15521 15853 15555
rect 15887 15521 15899 15555
rect 15841 15515 15899 15521
rect 14185 15487 14243 15493
rect 14185 15453 14197 15487
rect 14231 15453 14243 15487
rect 14185 15447 14243 15453
rect 14366 15444 14372 15496
rect 14424 15444 14430 15496
rect 14553 15487 14611 15493
rect 14553 15453 14565 15487
rect 14599 15484 14611 15487
rect 14642 15484 14648 15496
rect 14599 15456 14648 15484
rect 14599 15453 14611 15456
rect 14553 15447 14611 15453
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 15657 15487 15715 15493
rect 15657 15478 15669 15487
rect 15488 15453 15669 15478
rect 15703 15453 15715 15487
rect 15488 15450 15715 15453
rect 6362 15416 6368 15428
rect 6196 15388 6368 15416
rect 6362 15376 6368 15388
rect 6420 15376 6426 15428
rect 6454 15376 6460 15428
rect 6512 15376 6518 15428
rect 6914 15376 6920 15428
rect 6972 15376 6978 15428
rect 12161 15419 12219 15425
rect 7760 15388 11008 15416
rect 5442 15308 5448 15360
rect 5500 15348 5506 15360
rect 7760 15348 7788 15388
rect 10980 15357 11008 15388
rect 12161 15385 12173 15419
rect 12207 15416 12219 15419
rect 12434 15416 12440 15428
rect 12207 15388 12440 15416
rect 12207 15385 12219 15388
rect 12161 15379 12219 15385
rect 12434 15376 12440 15388
rect 12492 15376 12498 15428
rect 13909 15419 13967 15425
rect 12544 15388 12650 15416
rect 5500 15320 7788 15348
rect 10965 15351 11023 15357
rect 5500 15308 5506 15320
rect 10965 15317 10977 15351
rect 11011 15317 11023 15351
rect 10965 15311 11023 15317
rect 11425 15351 11483 15357
rect 11425 15317 11437 15351
rect 11471 15348 11483 15351
rect 11514 15348 11520 15360
rect 11471 15320 11520 15348
rect 11471 15317 11483 15320
rect 11425 15311 11483 15317
rect 11514 15308 11520 15320
rect 11572 15308 11578 15360
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 12250 15348 12256 15360
rect 11756 15320 12256 15348
rect 11756 15308 11762 15320
rect 12250 15308 12256 15320
rect 12308 15348 12314 15360
rect 12544 15348 12572 15388
rect 13909 15385 13921 15419
rect 13955 15416 13967 15419
rect 14384 15416 14412 15444
rect 13955 15388 14412 15416
rect 13955 15385 13967 15388
rect 13909 15379 13967 15385
rect 12308 15320 12572 15348
rect 15488 15348 15516 15450
rect 15657 15447 15715 15450
rect 15930 15444 15936 15496
rect 15988 15484 15994 15496
rect 16040 15484 16068 15592
rect 17678 15580 17684 15592
rect 17736 15580 17742 15632
rect 18874 15620 18880 15632
rect 17972 15592 18880 15620
rect 17972 15564 18000 15592
rect 18874 15580 18880 15592
rect 18932 15580 18938 15632
rect 18966 15580 18972 15632
rect 19024 15620 19030 15632
rect 19024 15592 19840 15620
rect 19024 15580 19030 15592
rect 16390 15512 16396 15564
rect 16448 15512 16454 15564
rect 16758 15512 16764 15564
rect 16816 15552 16822 15564
rect 16942 15552 16948 15564
rect 16816 15524 16948 15552
rect 16816 15512 16822 15524
rect 16942 15512 16948 15524
rect 17000 15512 17006 15564
rect 17954 15512 17960 15564
rect 18012 15512 18018 15564
rect 18598 15512 18604 15564
rect 18656 15552 18662 15564
rect 18785 15555 18843 15561
rect 18785 15552 18797 15555
rect 18656 15524 18797 15552
rect 18656 15512 18662 15524
rect 18785 15521 18797 15524
rect 18831 15521 18843 15555
rect 18785 15515 18843 15521
rect 18892 15524 19380 15552
rect 15988 15456 16068 15484
rect 16109 15489 16167 15495
rect 15988 15444 15994 15456
rect 16109 15455 16121 15489
rect 16155 15455 16167 15489
rect 16109 15449 16167 15455
rect 16301 15487 16359 15493
rect 16301 15453 16313 15487
rect 16347 15484 16359 15487
rect 16408 15484 16436 15512
rect 18892 15484 18920 15524
rect 19352 15493 19380 15524
rect 16347 15456 16436 15484
rect 18248 15456 18920 15484
rect 18969 15487 19027 15493
rect 16347 15453 16359 15456
rect 15746 15376 15752 15428
rect 15804 15416 15810 15428
rect 16132 15416 16160 15449
rect 16301 15447 16359 15453
rect 18248 15428 18276 15456
rect 18969 15453 18981 15487
rect 19015 15453 19027 15487
rect 18969 15447 19027 15453
rect 19061 15487 19119 15493
rect 19061 15453 19073 15487
rect 19107 15453 19119 15487
rect 19061 15447 19119 15453
rect 19337 15487 19395 15493
rect 19337 15453 19349 15487
rect 19383 15453 19395 15487
rect 19337 15447 19395 15453
rect 15804 15388 16160 15416
rect 15804 15376 15810 15388
rect 18230 15376 18236 15428
rect 18288 15376 18294 15428
rect 18417 15419 18475 15425
rect 18417 15385 18429 15419
rect 18463 15416 18475 15419
rect 18463 15388 18644 15416
rect 18463 15385 18475 15388
rect 18417 15379 18475 15385
rect 18616 15357 18644 15388
rect 18782 15376 18788 15428
rect 18840 15416 18846 15428
rect 18984 15416 19012 15447
rect 18840 15388 19012 15416
rect 19076 15416 19104 15447
rect 19426 15444 19432 15496
rect 19484 15444 19490 15496
rect 19812 15484 19840 15592
rect 23952 15592 24992 15620
rect 20809 15555 20867 15561
rect 20809 15521 20821 15555
rect 20855 15552 20867 15555
rect 21082 15552 21088 15564
rect 20855 15524 21088 15552
rect 20855 15521 20867 15524
rect 20809 15515 20867 15521
rect 21082 15512 21088 15524
rect 21140 15512 21146 15564
rect 22646 15512 22652 15564
rect 22704 15552 22710 15564
rect 22704 15524 23428 15552
rect 22704 15512 22710 15524
rect 19981 15487 20039 15493
rect 19981 15484 19993 15487
rect 19812 15456 19993 15484
rect 19981 15453 19993 15456
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 20717 15487 20775 15493
rect 20717 15453 20729 15487
rect 20763 15453 20775 15487
rect 20717 15447 20775 15453
rect 19444 15416 19472 15444
rect 20070 15416 20076 15428
rect 19076 15388 20076 15416
rect 18840 15376 18846 15388
rect 20070 15376 20076 15388
rect 20128 15376 20134 15428
rect 16117 15351 16175 15357
rect 16117 15348 16129 15351
rect 15488 15320 16129 15348
rect 12308 15308 12314 15320
rect 16117 15317 16129 15320
rect 16163 15317 16175 15351
rect 16117 15311 16175 15317
rect 18601 15351 18659 15357
rect 18601 15317 18613 15351
rect 18647 15348 18659 15351
rect 18966 15348 18972 15360
rect 18647 15320 18972 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 18966 15308 18972 15320
rect 19024 15308 19030 15360
rect 19334 15308 19340 15360
rect 19392 15308 19398 15360
rect 19978 15308 19984 15360
rect 20036 15348 20042 15360
rect 20530 15348 20536 15360
rect 20036 15320 20536 15348
rect 20036 15308 20042 15320
rect 20530 15308 20536 15320
rect 20588 15348 20594 15360
rect 20732 15348 20760 15447
rect 22002 15444 22008 15496
rect 22060 15484 22066 15496
rect 22925 15487 22983 15493
rect 22925 15484 22937 15487
rect 22060 15456 22937 15484
rect 22060 15444 22066 15456
rect 22925 15453 22937 15456
rect 22971 15453 22983 15487
rect 22925 15447 22983 15453
rect 23014 15444 23020 15496
rect 23072 15484 23078 15496
rect 23400 15493 23428 15524
rect 23952 15496 23980 15592
rect 23109 15487 23167 15493
rect 23109 15484 23121 15487
rect 23072 15456 23121 15484
rect 23072 15444 23078 15456
rect 23109 15453 23121 15456
rect 23155 15453 23167 15487
rect 23109 15447 23167 15453
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15453 23719 15487
rect 23661 15447 23719 15453
rect 23753 15487 23811 15493
rect 23753 15453 23765 15487
rect 23799 15484 23811 15487
rect 23934 15484 23940 15496
rect 23799 15456 23940 15484
rect 23799 15453 23811 15456
rect 23753 15447 23811 15453
rect 23676 15416 23704 15447
rect 23934 15444 23940 15456
rect 23992 15444 23998 15496
rect 24486 15444 24492 15496
rect 24544 15444 24550 15496
rect 24670 15444 24676 15496
rect 24728 15484 24734 15496
rect 24964 15493 24992 15592
rect 24765 15487 24823 15493
rect 24765 15484 24777 15487
rect 24728 15456 24777 15484
rect 24728 15444 24734 15456
rect 24765 15453 24777 15456
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 24949 15487 25007 15493
rect 24949 15453 24961 15487
rect 24995 15484 25007 15487
rect 25222 15484 25228 15496
rect 24995 15456 25228 15484
rect 24995 15453 25007 15456
rect 24949 15447 25007 15453
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 25424 15493 25452 15660
rect 26329 15657 26341 15691
rect 26375 15688 26387 15691
rect 27338 15688 27344 15700
rect 26375 15660 27344 15688
rect 26375 15657 26387 15660
rect 26329 15651 26387 15657
rect 27338 15648 27344 15660
rect 27396 15648 27402 15700
rect 29454 15648 29460 15700
rect 29512 15648 29518 15700
rect 30742 15648 30748 15700
rect 30800 15648 30806 15700
rect 31386 15648 31392 15700
rect 31444 15648 31450 15700
rect 32214 15648 32220 15700
rect 32272 15688 32278 15700
rect 32309 15691 32367 15697
rect 32309 15688 32321 15691
rect 32272 15660 32321 15688
rect 32272 15648 32278 15660
rect 32309 15657 32321 15660
rect 32355 15657 32367 15691
rect 32309 15651 32367 15657
rect 32582 15648 32588 15700
rect 32640 15688 32646 15700
rect 32769 15691 32827 15697
rect 32769 15688 32781 15691
rect 32640 15660 32781 15688
rect 32640 15648 32646 15660
rect 32769 15657 32781 15660
rect 32815 15657 32827 15691
rect 32769 15651 32827 15657
rect 32858 15648 32864 15700
rect 32916 15688 32922 15700
rect 33229 15691 33287 15697
rect 33229 15688 33241 15691
rect 32916 15660 33241 15688
rect 32916 15648 32922 15660
rect 33229 15657 33241 15660
rect 33275 15657 33287 15691
rect 33229 15651 33287 15657
rect 34790 15648 34796 15700
rect 34848 15688 34854 15700
rect 35161 15691 35219 15697
rect 35161 15688 35173 15691
rect 34848 15660 35173 15688
rect 34848 15648 34854 15660
rect 35161 15657 35173 15660
rect 35207 15657 35219 15691
rect 35161 15651 35219 15657
rect 35437 15691 35495 15697
rect 35437 15657 35449 15691
rect 35483 15688 35495 15691
rect 35526 15688 35532 15700
rect 35483 15660 35532 15688
rect 35483 15657 35495 15660
rect 35437 15651 35495 15657
rect 35526 15648 35532 15660
rect 35584 15648 35590 15700
rect 26605 15623 26663 15629
rect 26605 15589 26617 15623
rect 26651 15620 26663 15623
rect 26651 15592 27108 15620
rect 26651 15589 26663 15592
rect 26605 15583 26663 15589
rect 27080 15496 27108 15592
rect 27172 15592 28764 15620
rect 27172 15564 27200 15592
rect 27154 15512 27160 15564
rect 27212 15512 27218 15564
rect 27430 15512 27436 15564
rect 27488 15552 27494 15564
rect 27709 15555 27767 15561
rect 27488 15524 27660 15552
rect 27488 15512 27494 15524
rect 25409 15487 25467 15493
rect 25409 15453 25421 15487
rect 25455 15453 25467 15487
rect 25409 15447 25467 15453
rect 25498 15444 25504 15496
rect 25556 15484 25562 15496
rect 25961 15487 26019 15493
rect 25961 15484 25973 15487
rect 25556 15456 25973 15484
rect 25556 15444 25562 15456
rect 25961 15453 25973 15456
rect 26007 15453 26019 15487
rect 25961 15447 26019 15453
rect 26050 15444 26056 15496
rect 26108 15484 26114 15496
rect 26145 15487 26203 15493
rect 26145 15484 26157 15487
rect 26108 15456 26157 15484
rect 26108 15444 26114 15456
rect 26145 15453 26157 15456
rect 26191 15453 26203 15487
rect 26145 15447 26203 15453
rect 26234 15444 26240 15496
rect 26292 15484 26298 15496
rect 26421 15487 26479 15493
rect 26421 15484 26433 15487
rect 26292 15456 26433 15484
rect 26292 15444 26298 15456
rect 26421 15453 26433 15456
rect 26467 15453 26479 15487
rect 26421 15447 26479 15453
rect 27062 15444 27068 15496
rect 27120 15484 27126 15496
rect 27632 15493 27660 15524
rect 27709 15521 27721 15555
rect 27755 15552 27767 15555
rect 27985 15555 28043 15561
rect 27985 15552 27997 15555
rect 27755 15524 27997 15552
rect 27755 15521 27767 15524
rect 27709 15515 27767 15521
rect 27985 15521 27997 15524
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 27617 15487 27675 15493
rect 27120 15456 27568 15484
rect 27120 15444 27126 15456
rect 27430 15416 27436 15428
rect 23676 15388 27436 15416
rect 27430 15376 27436 15388
rect 27488 15376 27494 15428
rect 20588 15320 20760 15348
rect 20588 15308 20594 15320
rect 24670 15308 24676 15360
rect 24728 15348 24734 15360
rect 25498 15348 25504 15360
rect 24728 15320 25504 15348
rect 24728 15308 24734 15320
rect 25498 15308 25504 15320
rect 25556 15308 25562 15360
rect 25593 15351 25651 15357
rect 25593 15317 25605 15351
rect 25639 15348 25651 15351
rect 25682 15348 25688 15360
rect 25639 15320 25688 15348
rect 25639 15317 25651 15320
rect 25593 15311 25651 15317
rect 25682 15308 25688 15320
rect 25740 15308 25746 15360
rect 27249 15351 27307 15357
rect 27249 15317 27261 15351
rect 27295 15348 27307 15351
rect 27338 15348 27344 15360
rect 27295 15320 27344 15348
rect 27295 15317 27307 15320
rect 27249 15311 27307 15317
rect 27338 15308 27344 15320
rect 27396 15308 27402 15360
rect 27540 15348 27568 15456
rect 27617 15453 27629 15487
rect 27663 15484 27675 15487
rect 28074 15484 28080 15496
rect 27663 15456 28080 15484
rect 27663 15453 27675 15456
rect 27617 15447 27675 15453
rect 28074 15444 28080 15456
rect 28132 15444 28138 15496
rect 28736 15493 28764 15592
rect 29472 15552 29500 15648
rect 29472 15524 29868 15552
rect 28169 15487 28227 15493
rect 28169 15453 28181 15487
rect 28215 15453 28227 15487
rect 28169 15447 28227 15453
rect 28445 15487 28503 15493
rect 28445 15453 28457 15487
rect 28491 15484 28503 15487
rect 28629 15487 28687 15493
rect 28629 15484 28641 15487
rect 28491 15456 28641 15484
rect 28491 15453 28503 15456
rect 28445 15447 28503 15453
rect 28629 15453 28641 15456
rect 28675 15453 28687 15487
rect 28629 15447 28687 15453
rect 28721 15487 28779 15493
rect 28721 15453 28733 15487
rect 28767 15484 28779 15487
rect 29086 15484 29092 15496
rect 28767 15456 29092 15484
rect 28767 15453 28779 15456
rect 28721 15447 28779 15453
rect 28184 15416 28212 15447
rect 29086 15444 29092 15456
rect 29144 15484 29150 15496
rect 29840 15493 29868 15524
rect 29641 15487 29699 15493
rect 29641 15484 29653 15487
rect 29144 15456 29653 15484
rect 29144 15444 29150 15456
rect 29641 15453 29653 15456
rect 29687 15453 29699 15487
rect 29641 15447 29699 15453
rect 29825 15487 29883 15493
rect 29825 15453 29837 15487
rect 29871 15453 29883 15487
rect 30760 15484 30788 15648
rect 31404 15552 31432 15648
rect 32401 15623 32459 15629
rect 32401 15589 32413 15623
rect 32447 15620 32459 15623
rect 32447 15592 33456 15620
rect 32447 15589 32459 15592
rect 32401 15583 32459 15589
rect 31849 15555 31907 15561
rect 31404 15524 31708 15552
rect 31680 15493 31708 15524
rect 31849 15521 31861 15555
rect 31895 15552 31907 15555
rect 32217 15555 32275 15561
rect 32217 15552 32229 15555
rect 31895 15524 32229 15552
rect 31895 15521 31907 15524
rect 31849 15515 31907 15521
rect 32217 15521 32229 15524
rect 32263 15552 32275 15555
rect 33321 15555 33379 15561
rect 33321 15552 33333 15555
rect 32263 15524 33333 15552
rect 32263 15521 32275 15524
rect 32217 15515 32275 15521
rect 33321 15521 33333 15524
rect 33367 15521 33379 15555
rect 33321 15515 33379 15521
rect 33428 15496 33456 15592
rect 34790 15512 34796 15564
rect 34848 15512 34854 15564
rect 35618 15512 35624 15564
rect 35676 15512 35682 15564
rect 31481 15487 31539 15493
rect 31481 15484 31493 15487
rect 30760 15456 31493 15484
rect 29825 15447 29883 15453
rect 31481 15453 31493 15456
rect 31527 15453 31539 15487
rect 31481 15447 31539 15453
rect 31665 15487 31723 15493
rect 31665 15453 31677 15487
rect 31711 15453 31723 15487
rect 31665 15447 31723 15453
rect 32493 15487 32551 15493
rect 32493 15453 32505 15487
rect 32539 15484 32551 15487
rect 32858 15484 32864 15496
rect 32539 15456 32864 15484
rect 32539 15453 32551 15456
rect 32493 15447 32551 15453
rect 32858 15444 32864 15456
rect 32916 15444 32922 15496
rect 33410 15444 33416 15496
rect 33468 15444 33474 15496
rect 34606 15444 34612 15496
rect 34664 15444 34670 15496
rect 34698 15444 34704 15496
rect 34756 15484 34762 15496
rect 34885 15487 34943 15493
rect 34885 15484 34897 15487
rect 34756 15456 34897 15484
rect 34756 15444 34762 15456
rect 34885 15453 34897 15456
rect 34931 15453 34943 15487
rect 34885 15447 34943 15453
rect 35713 15487 35771 15493
rect 35713 15453 35725 15487
rect 35759 15453 35771 15487
rect 35713 15447 35771 15453
rect 30282 15416 30288 15428
rect 28184 15388 30288 15416
rect 30282 15376 30288 15388
rect 30340 15376 30346 15428
rect 32214 15376 32220 15428
rect 32272 15416 32278 15428
rect 32737 15419 32795 15425
rect 32737 15416 32749 15419
rect 32272 15388 32749 15416
rect 32272 15376 32278 15388
rect 32737 15385 32749 15388
rect 32783 15385 32795 15419
rect 32737 15379 32795 15385
rect 32953 15419 33011 15425
rect 32953 15385 32965 15419
rect 32999 15416 33011 15419
rect 34624 15416 34652 15444
rect 35728 15416 35756 15447
rect 32999 15388 33088 15416
rect 34624 15388 35756 15416
rect 32999 15385 33011 15388
rect 32953 15379 33011 15385
rect 28350 15348 28356 15360
rect 27540 15320 28356 15348
rect 28350 15308 28356 15320
rect 28408 15308 28414 15360
rect 30650 15308 30656 15360
rect 30708 15308 30714 15360
rect 32582 15308 32588 15360
rect 32640 15308 32646 15360
rect 33060 15357 33088 15388
rect 33045 15351 33103 15357
rect 33045 15317 33057 15351
rect 33091 15317 33103 15351
rect 33045 15311 33103 15317
rect 1104 15258 38272 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38272 15258
rect 1104 15184 38272 15206
rect 2961 15147 3019 15153
rect 2961 15113 2973 15147
rect 3007 15144 3019 15147
rect 3697 15147 3755 15153
rect 3697 15144 3709 15147
rect 3007 15116 3709 15144
rect 3007 15113 3019 15116
rect 2961 15107 3019 15113
rect 3697 15113 3709 15116
rect 3743 15113 3755 15147
rect 3697 15107 3755 15113
rect 4065 15147 4123 15153
rect 4065 15113 4077 15147
rect 4111 15144 4123 15147
rect 5442 15144 5448 15156
rect 4111 15116 5448 15144
rect 4111 15113 4123 15116
rect 4065 15107 4123 15113
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 6454 15104 6460 15156
rect 6512 15144 6518 15156
rect 6641 15147 6699 15153
rect 6641 15144 6653 15147
rect 6512 15116 6653 15144
rect 6512 15104 6518 15116
rect 6641 15113 6653 15116
rect 6687 15113 6699 15147
rect 6641 15107 6699 15113
rect 7558 15104 7564 15156
rect 7616 15104 7622 15156
rect 8294 15104 8300 15156
rect 8352 15104 8358 15156
rect 8754 15104 8760 15156
rect 8812 15104 8818 15156
rect 9490 15104 9496 15156
rect 9548 15104 9554 15156
rect 11977 15147 12035 15153
rect 11977 15113 11989 15147
rect 12023 15144 12035 15147
rect 12158 15144 12164 15156
rect 12023 15116 12164 15144
rect 12023 15113 12035 15116
rect 11977 15107 12035 15113
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 13909 15147 13967 15153
rect 13909 15144 13921 15147
rect 12492 15116 13921 15144
rect 12492 15104 12498 15116
rect 13909 15113 13921 15116
rect 13955 15113 13967 15147
rect 13909 15107 13967 15113
rect 14550 15104 14556 15156
rect 14608 15144 14614 15156
rect 14918 15144 14924 15156
rect 14608 15116 14924 15144
rect 14608 15104 14614 15116
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 15749 15147 15807 15153
rect 15749 15113 15761 15147
rect 15795 15144 15807 15147
rect 16390 15144 16396 15156
rect 15795 15116 16396 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 18782 15104 18788 15156
rect 18840 15104 18846 15156
rect 26050 15104 26056 15156
rect 26108 15104 26114 15156
rect 27065 15147 27123 15153
rect 27065 15113 27077 15147
rect 27111 15144 27123 15147
rect 27338 15144 27344 15156
rect 27111 15116 27344 15144
rect 27111 15113 27123 15116
rect 27065 15107 27123 15113
rect 27338 15104 27344 15116
rect 27396 15144 27402 15156
rect 27614 15144 27620 15156
rect 27396 15116 27620 15144
rect 27396 15104 27402 15116
rect 27614 15104 27620 15116
rect 27672 15104 27678 15156
rect 27890 15104 27896 15156
rect 27948 15144 27954 15156
rect 32582 15144 32588 15156
rect 27948 15116 32588 15144
rect 27948 15104 27954 15116
rect 32582 15104 32588 15116
rect 32640 15104 32646 15156
rect 34333 15147 34391 15153
rect 34333 15113 34345 15147
rect 34379 15144 34391 15147
rect 34790 15144 34796 15156
rect 34379 15116 34796 15144
rect 34379 15113 34391 15116
rect 34333 15107 34391 15113
rect 34790 15104 34796 15116
rect 34848 15104 34854 15156
rect 4154 15076 4160 15088
rect 3436 15048 4160 15076
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 15008 2927 15011
rect 3234 15008 3240 15020
rect 2915 14980 3240 15008
rect 2915 14977 2927 14980
rect 2869 14971 2927 14977
rect 3234 14968 3240 14980
rect 3292 15008 3298 15020
rect 3436 15017 3464 15048
rect 4154 15036 4160 15048
rect 4212 15076 4218 15088
rect 4212 15048 4568 15076
rect 4212 15036 4218 15048
rect 3421 15011 3479 15017
rect 3421 15008 3433 15011
rect 3292 14980 3433 15008
rect 3292 14968 3298 14980
rect 3421 14977 3433 14980
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 15008 3663 15011
rect 3970 15008 3976 15020
rect 3651 14980 3976 15008
rect 3651 14977 3663 14980
rect 3605 14971 3663 14977
rect 3970 14968 3976 14980
rect 4028 15008 4034 15020
rect 4028 14980 4384 15008
rect 4028 14968 4034 14980
rect 3142 14900 3148 14952
rect 3200 14900 3206 14952
rect 4157 14943 4215 14949
rect 4157 14940 4169 14943
rect 4080 14912 4169 14940
rect 4080 14884 4108 14912
rect 4157 14909 4169 14912
rect 4203 14909 4215 14943
rect 4157 14903 4215 14909
rect 4246 14900 4252 14952
rect 4304 14900 4310 14952
rect 4062 14832 4068 14884
rect 4120 14832 4126 14884
rect 2498 14764 2504 14816
rect 2556 14764 2562 14816
rect 3602 14764 3608 14816
rect 3660 14764 3666 14816
rect 3878 14764 3884 14816
rect 3936 14804 3942 14816
rect 4264 14804 4292 14900
rect 4356 14872 4384 14980
rect 4540 14949 4568 15048
rect 4614 15036 4620 15088
rect 4672 15076 4678 15088
rect 4893 15079 4951 15085
rect 4893 15076 4905 15079
rect 4672 15048 4905 15076
rect 4672 15036 4678 15048
rect 4893 15045 4905 15048
rect 4939 15045 4951 15079
rect 4893 15039 4951 15045
rect 4706 14968 4712 15020
rect 4764 14968 4770 15020
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 7469 15011 7527 15017
rect 6871 14980 7144 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14909 4583 14943
rect 4525 14903 4583 14909
rect 4724 14872 4752 14968
rect 7116 14881 7144 14980
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 8113 15011 8171 15017
rect 7515 14980 8064 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 7190 14900 7196 14952
rect 7248 14940 7254 14952
rect 7653 14943 7711 14949
rect 7653 14940 7665 14943
rect 7248 14912 7665 14940
rect 7248 14900 7254 14912
rect 7653 14909 7665 14912
rect 7699 14909 7711 14943
rect 7653 14903 7711 14909
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14909 7987 14943
rect 8036 14940 8064 14980
rect 8113 14977 8125 15011
rect 8159 15008 8171 15011
rect 8312 15008 8340 15104
rect 8159 14980 8340 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8386 14968 8392 15020
rect 8444 15008 8450 15020
rect 8772 15008 8800 15104
rect 9033 15079 9091 15085
rect 9033 15076 9045 15079
rect 8956 15048 9045 15076
rect 8956 15020 8984 15048
rect 9033 15045 9045 15048
rect 9079 15045 9091 15079
rect 9033 15039 9091 15045
rect 8444 14980 8800 15008
rect 8444 14968 8450 14980
rect 8938 14968 8944 15020
rect 8996 14968 9002 15020
rect 9508 15008 9536 15104
rect 9582 15036 9588 15088
rect 9640 15076 9646 15088
rect 10778 15076 10784 15088
rect 9640 15048 10784 15076
rect 9640 15036 9646 15048
rect 10778 15036 10784 15048
rect 10836 15076 10842 15088
rect 11885 15079 11943 15085
rect 11885 15076 11897 15079
rect 10836 15048 11897 15076
rect 10836 15036 10842 15048
rect 11885 15045 11897 15048
rect 11931 15045 11943 15079
rect 14568 15076 14596 15104
rect 11885 15039 11943 15045
rect 13004 15048 13768 15076
rect 13004 15017 13032 15048
rect 13740 15020 13768 15048
rect 13832 15048 14228 15076
rect 13832 15020 13860 15048
rect 10505 15011 10563 15017
rect 9508 14980 9628 15008
rect 8297 14943 8355 14949
rect 8297 14940 8309 14943
rect 8036 14912 8309 14940
rect 7929 14903 7987 14909
rect 8297 14909 8309 14912
rect 8343 14940 8355 14943
rect 9490 14940 9496 14952
rect 8343 14912 9496 14940
rect 8343 14909 8355 14912
rect 8297 14903 8355 14909
rect 4356 14844 4752 14872
rect 7101 14875 7159 14881
rect 7101 14841 7113 14875
rect 7147 14841 7159 14875
rect 7944 14872 7972 14903
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 9600 14949 9628 14980
rect 10505 14977 10517 15011
rect 10551 15008 10563 15011
rect 12989 15011 13047 15017
rect 10551 14980 11560 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 9585 14943 9643 14949
rect 9585 14909 9597 14943
rect 9631 14909 9643 14943
rect 9585 14903 9643 14909
rect 8110 14872 8116 14884
rect 7944 14844 8116 14872
rect 7101 14835 7159 14841
rect 8110 14832 8116 14844
rect 8168 14832 8174 14884
rect 9030 14832 9036 14884
rect 9088 14832 9094 14884
rect 11532 14881 11560 14980
rect 12989 14977 13001 15011
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 13354 14968 13360 15020
rect 13412 14968 13418 15020
rect 13722 14968 13728 15020
rect 13780 14968 13786 15020
rect 13814 14968 13820 15020
rect 13872 14968 13878 15020
rect 14090 14968 14096 15020
rect 14148 14968 14154 15020
rect 14200 15017 14228 15048
rect 14292 15048 14596 15076
rect 14737 15079 14795 15085
rect 14292 15017 14320 15048
rect 14737 15045 14749 15079
rect 14783 15076 14795 15079
rect 15013 15079 15071 15085
rect 15013 15076 15025 15079
rect 14783 15048 15025 15076
rect 14783 15045 14795 15048
rect 14737 15039 14795 15045
rect 15013 15045 15025 15048
rect 15059 15045 15071 15079
rect 15013 15039 15071 15045
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 14461 15011 14519 15017
rect 14461 15008 14473 15011
rect 14424 14980 14473 15008
rect 14424 14968 14430 14980
rect 14461 14977 14473 14980
rect 14507 14977 14519 15011
rect 14461 14971 14519 14977
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 14829 15011 14887 15017
rect 14829 14977 14841 15011
rect 14875 15008 14887 15011
rect 15105 15011 15163 15017
rect 14875 14980 14964 15008
rect 14875 14977 14887 14980
rect 14829 14971 14887 14977
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 12618 14940 12624 14952
rect 12207 14912 12624 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 12618 14900 12624 14912
rect 12676 14900 12682 14952
rect 12802 14900 12808 14952
rect 12860 14940 12866 14952
rect 14568 14940 14596 14971
rect 12860 14912 14596 14940
rect 12860 14900 12866 14912
rect 14292 14884 14320 14912
rect 14642 14900 14648 14952
rect 14700 14940 14706 14952
rect 14936 14940 14964 14980
rect 15105 14977 15117 15011
rect 15151 14977 15163 15011
rect 15105 14971 15163 14977
rect 15010 14940 15016 14952
rect 14700 14912 14872 14940
rect 14936 14912 15016 14940
rect 14700 14900 14706 14912
rect 11517 14875 11575 14881
rect 11517 14841 11529 14875
rect 11563 14841 11575 14875
rect 11517 14835 11575 14841
rect 14274 14832 14280 14884
rect 14332 14832 14338 14884
rect 14844 14881 14872 14912
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 14829 14875 14887 14881
rect 14829 14841 14841 14875
rect 14875 14841 14887 14875
rect 15120 14872 15148 14971
rect 15470 14968 15476 15020
rect 15528 14968 15534 15020
rect 15565 15011 15623 15017
rect 15565 14977 15577 15011
rect 15611 15008 15623 15011
rect 15930 15008 15936 15020
rect 15611 14980 15936 15008
rect 15611 14977 15623 14980
rect 15565 14971 15623 14977
rect 15930 14968 15936 14980
rect 15988 15008 15994 15020
rect 16114 15008 16120 15020
rect 15988 14980 16120 15008
rect 15988 14968 15994 14980
rect 16114 14968 16120 14980
rect 16172 14968 16178 15020
rect 16206 14968 16212 15020
rect 16264 14968 16270 15020
rect 16408 15008 16436 15104
rect 18800 15076 18828 15104
rect 20438 15076 20444 15088
rect 16960 15048 19196 15076
rect 16960 15020 16988 15048
rect 16485 15011 16543 15017
rect 16485 15008 16497 15011
rect 16408 14980 16497 15008
rect 16485 14977 16497 14980
rect 16531 14977 16543 15011
rect 16485 14971 16543 14977
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 15008 16911 15011
rect 16942 15008 16948 15020
rect 16899 14980 16948 15008
rect 16899 14977 16911 14980
rect 16853 14971 16911 14977
rect 16942 14968 16948 14980
rect 17000 14968 17006 15020
rect 17034 14968 17040 15020
rect 17092 14968 17098 15020
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 14977 17187 15011
rect 17129 14971 17187 14977
rect 16298 14900 16304 14952
rect 16356 14940 16362 14952
rect 17144 14940 17172 14971
rect 17218 14968 17224 15020
rect 17276 15008 17282 15020
rect 17405 15011 17463 15017
rect 17405 15008 17417 15011
rect 17276 14980 17417 15008
rect 17276 14968 17282 14980
rect 17405 14977 17417 14980
rect 17451 14977 17463 15011
rect 17405 14971 17463 14977
rect 17678 14968 17684 15020
rect 17736 14968 17742 15020
rect 18598 14968 18604 15020
rect 18656 15008 18662 15020
rect 19168 15017 19196 15048
rect 20180 15048 20444 15076
rect 20180 15020 20208 15048
rect 20438 15036 20444 15048
rect 20496 15036 20502 15088
rect 26068 15076 26096 15104
rect 28997 15079 29055 15085
rect 25516 15048 26096 15076
rect 18785 15011 18843 15017
rect 18785 15008 18797 15011
rect 18656 14980 18797 15008
rect 18656 14968 18662 14980
rect 18785 14977 18797 14980
rect 18831 14977 18843 15011
rect 18785 14971 18843 14977
rect 19153 15011 19211 15017
rect 19153 14977 19165 15011
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19521 15011 19579 15017
rect 19521 15008 19533 15011
rect 19484 14980 19533 15008
rect 19484 14968 19490 14980
rect 19521 14977 19533 14980
rect 19567 14977 19579 15011
rect 19521 14971 19579 14977
rect 19978 14968 19984 15020
rect 20036 15008 20042 15020
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 20036 14980 20085 15008
rect 20036 14968 20042 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20162 14968 20168 15020
rect 20220 14968 20226 15020
rect 20349 15011 20407 15017
rect 20349 14977 20361 15011
rect 20395 15008 20407 15011
rect 20806 15008 20812 15020
rect 20395 14980 20812 15008
rect 20395 14977 20407 14980
rect 20349 14971 20407 14977
rect 16356 14912 17172 14940
rect 18141 14943 18199 14949
rect 16356 14900 16362 14912
rect 18141 14909 18153 14943
rect 18187 14940 18199 14943
rect 18230 14940 18236 14952
rect 18187 14912 18236 14940
rect 18187 14909 18199 14912
rect 18141 14903 18199 14909
rect 18230 14900 18236 14912
rect 18288 14900 18294 14952
rect 20364 14940 20392 14971
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 15008 22063 15011
rect 22189 15011 22247 15017
rect 22051 14980 22140 15008
rect 22051 14977 22063 14980
rect 22005 14971 22063 14977
rect 22112 14952 22140 14980
rect 22189 14977 22201 15011
rect 22235 15008 22247 15011
rect 22649 15011 22707 15017
rect 22649 15008 22661 15011
rect 22235 14980 22661 15008
rect 22235 14977 22247 14980
rect 22189 14971 22247 14977
rect 22649 14977 22661 14980
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 23198 14968 23204 15020
rect 23256 14968 23262 15020
rect 25516 15017 25544 15048
rect 25501 15011 25559 15017
rect 25501 14977 25513 15011
rect 25547 14977 25559 15011
rect 25501 14971 25559 14977
rect 25682 14968 25688 15020
rect 25740 15008 25746 15020
rect 25777 15011 25835 15017
rect 25777 15008 25789 15011
rect 25740 14980 25789 15008
rect 25740 14968 25746 14980
rect 25777 14977 25789 14980
rect 25823 14977 25835 15011
rect 25777 14971 25835 14977
rect 25961 15011 26019 15017
rect 25961 14977 25973 15011
rect 26007 15008 26019 15011
rect 26068 15008 26096 15048
rect 28552 15048 28948 15076
rect 26007 14980 26096 15008
rect 26007 14977 26019 14980
rect 25961 14971 26019 14977
rect 18708 14912 20392 14940
rect 15933 14875 15991 14881
rect 15933 14872 15945 14875
rect 15120 14844 15945 14872
rect 14829 14835 14887 14841
rect 15933 14841 15945 14844
rect 15979 14841 15991 14875
rect 18708 14872 18736 14912
rect 21818 14900 21824 14952
rect 21876 14900 21882 14952
rect 22094 14900 22100 14952
rect 22152 14900 22158 14952
rect 25792 14940 25820 14971
rect 26326 14968 26332 15020
rect 26384 14968 26390 15020
rect 26418 14968 26424 15020
rect 26476 15008 26482 15020
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26476 14980 26985 15008
rect 26476 14968 26482 14980
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 26973 14971 27031 14977
rect 27154 14968 27160 15020
rect 27212 15008 27218 15020
rect 27249 15011 27307 15017
rect 27249 15008 27261 15011
rect 27212 14980 27261 15008
rect 27212 14968 27218 14980
rect 27249 14977 27261 14980
rect 27295 14977 27307 15011
rect 27249 14971 27307 14977
rect 27798 14968 27804 15020
rect 27856 14968 27862 15020
rect 28077 15011 28135 15017
rect 28077 14977 28089 15011
rect 28123 15008 28135 15011
rect 28261 15011 28319 15017
rect 28261 15008 28273 15011
rect 28123 14980 28273 15008
rect 28123 14977 28135 14980
rect 28077 14971 28135 14977
rect 28261 14977 28273 14980
rect 28307 14977 28319 15011
rect 28261 14971 28319 14977
rect 26142 14940 26148 14952
rect 25792 14912 26148 14940
rect 26142 14900 26148 14912
rect 26200 14940 26206 14952
rect 26344 14940 26372 14968
rect 26200 14912 26372 14940
rect 27897 14943 27955 14949
rect 26200 14900 26206 14912
rect 27897 14909 27909 14943
rect 27943 14940 27955 14943
rect 28166 14940 28172 14952
rect 27943 14912 28172 14940
rect 27943 14909 27955 14912
rect 27897 14903 27955 14909
rect 28166 14900 28172 14912
rect 28224 14900 28230 14952
rect 28276 14940 28304 14971
rect 28442 14968 28448 15020
rect 28500 14968 28506 15020
rect 28552 15017 28580 15048
rect 28537 15011 28595 15017
rect 28537 14977 28549 15011
rect 28583 14977 28595 15011
rect 28537 14971 28595 14977
rect 28629 15011 28687 15017
rect 28629 14977 28641 15011
rect 28675 15008 28687 15011
rect 28718 15008 28724 15020
rect 28675 14980 28724 15008
rect 28675 14977 28687 14980
rect 28629 14971 28687 14977
rect 28718 14968 28724 14980
rect 28776 14968 28782 15020
rect 28813 15011 28871 15017
rect 28813 14977 28825 15011
rect 28859 14977 28871 15011
rect 28920 15008 28948 15048
rect 28997 15045 29009 15079
rect 29043 15076 29055 15079
rect 29043 15048 34008 15076
rect 29043 15045 29055 15048
rect 28997 15039 29055 15045
rect 28920 14980 29960 15008
rect 28813 14971 28871 14977
rect 28276 14912 28488 14940
rect 28460 14884 28488 14912
rect 15933 14835 15991 14841
rect 16316 14844 18736 14872
rect 3936 14776 4292 14804
rect 3936 14764 3942 14776
rect 8662 14764 8668 14816
rect 8720 14764 8726 14816
rect 8849 14807 8907 14813
rect 8849 14773 8861 14807
rect 8895 14804 8907 14807
rect 8938 14804 8944 14816
rect 8895 14776 8944 14804
rect 8895 14773 8907 14776
rect 8849 14767 8907 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 9766 14764 9772 14816
rect 9824 14764 9830 14816
rect 10226 14764 10232 14816
rect 10284 14804 10290 14816
rect 10321 14807 10379 14813
rect 10321 14804 10333 14807
rect 10284 14776 10333 14804
rect 10284 14764 10290 14776
rect 10321 14773 10333 14776
rect 10367 14773 10379 14807
rect 10321 14767 10379 14773
rect 11974 14764 11980 14816
rect 12032 14804 12038 14816
rect 12529 14807 12587 14813
rect 12529 14804 12541 14807
rect 12032 14776 12541 14804
rect 12032 14764 12038 14776
rect 12529 14773 12541 14776
rect 12575 14804 12587 14807
rect 16316 14804 16344 14844
rect 18782 14832 18788 14884
rect 18840 14832 18846 14884
rect 19426 14832 19432 14884
rect 19484 14872 19490 14884
rect 24118 14872 24124 14884
rect 19484 14844 24124 14872
rect 19484 14832 19490 14844
rect 24118 14832 24124 14844
rect 24176 14832 24182 14884
rect 24762 14832 24768 14884
rect 24820 14872 24826 14884
rect 27433 14875 27491 14881
rect 24820 14844 26464 14872
rect 24820 14832 24826 14844
rect 12575 14776 16344 14804
rect 12575 14773 12587 14776
rect 12529 14767 12587 14773
rect 16390 14764 16396 14816
rect 16448 14804 16454 14816
rect 17678 14804 17684 14816
rect 16448 14776 17684 14804
rect 16448 14764 16454 14776
rect 17678 14764 17684 14776
rect 17736 14764 17742 14816
rect 20530 14764 20536 14816
rect 20588 14764 20594 14816
rect 20806 14764 20812 14816
rect 20864 14804 20870 14816
rect 22186 14804 22192 14816
rect 20864 14776 22192 14804
rect 20864 14764 20870 14776
rect 22186 14764 22192 14776
rect 22244 14764 22250 14816
rect 22278 14764 22284 14816
rect 22336 14804 22342 14816
rect 24578 14804 24584 14816
rect 22336 14776 24584 14804
rect 22336 14764 22342 14776
rect 24578 14764 24584 14776
rect 24636 14764 24642 14816
rect 25590 14764 25596 14816
rect 25648 14764 25654 14816
rect 25961 14807 26019 14813
rect 25961 14773 25973 14807
rect 26007 14804 26019 14807
rect 26326 14804 26332 14816
rect 26007 14776 26332 14804
rect 26007 14773 26019 14776
rect 25961 14767 26019 14773
rect 26326 14764 26332 14776
rect 26384 14764 26390 14816
rect 26436 14804 26464 14844
rect 27433 14841 27445 14875
rect 27479 14872 27491 14875
rect 27985 14875 28043 14881
rect 27479 14844 27844 14872
rect 27479 14841 27491 14844
rect 27433 14835 27491 14841
rect 27617 14807 27675 14813
rect 27617 14804 27629 14807
rect 26436 14776 27629 14804
rect 27617 14773 27629 14776
rect 27663 14773 27675 14807
rect 27816 14804 27844 14844
rect 27985 14841 27997 14875
rect 28031 14841 28043 14875
rect 27985 14835 28043 14841
rect 28000 14804 28028 14835
rect 28442 14832 28448 14884
rect 28500 14832 28506 14884
rect 28534 14832 28540 14884
rect 28592 14872 28598 14884
rect 28828 14872 28856 14971
rect 29932 14952 29960 14980
rect 30650 14968 30656 15020
rect 30708 14968 30714 15020
rect 30834 14968 30840 15020
rect 30892 14968 30898 15020
rect 30929 15011 30987 15017
rect 30929 14977 30941 15011
rect 30975 14977 30987 15011
rect 30929 14971 30987 14977
rect 29914 14900 29920 14952
rect 29972 14900 29978 14952
rect 30558 14900 30564 14952
rect 30616 14940 30622 14952
rect 30944 14940 30972 14971
rect 31110 14968 31116 15020
rect 31168 14968 31174 15020
rect 33042 14968 33048 15020
rect 33100 14968 33106 15020
rect 33980 15017 34008 15048
rect 33965 15011 34023 15017
rect 33965 14977 33977 15011
rect 34011 14977 34023 15011
rect 33965 14971 34023 14977
rect 30616 14912 30972 14940
rect 30616 14900 30622 14912
rect 32950 14900 32956 14952
rect 33008 14900 33014 14952
rect 33873 14943 33931 14949
rect 33873 14940 33885 14943
rect 33428 14912 33885 14940
rect 28592 14844 28856 14872
rect 28592 14832 28598 14844
rect 30466 14832 30472 14884
rect 30524 14872 30530 14884
rect 30742 14872 30748 14884
rect 30524 14844 30748 14872
rect 30524 14832 30530 14844
rect 30742 14832 30748 14844
rect 30800 14872 30806 14884
rect 33428 14881 33456 14912
rect 33873 14909 33885 14912
rect 33919 14909 33931 14943
rect 33873 14903 33931 14909
rect 30837 14875 30895 14881
rect 30837 14872 30849 14875
rect 30800 14844 30849 14872
rect 30800 14832 30806 14844
rect 30837 14841 30849 14844
rect 30883 14841 30895 14875
rect 33413 14875 33471 14881
rect 30837 14835 30895 14841
rect 30944 14844 31432 14872
rect 27816 14776 28028 14804
rect 27617 14767 27675 14773
rect 28810 14764 28816 14816
rect 28868 14804 28874 14816
rect 30944 14804 30972 14844
rect 31404 14816 31432 14844
rect 33413 14841 33425 14875
rect 33459 14841 33471 14875
rect 33413 14835 33471 14841
rect 28868 14776 30972 14804
rect 28868 14764 28874 14776
rect 31018 14764 31024 14816
rect 31076 14764 31082 14816
rect 31386 14764 31392 14816
rect 31444 14764 31450 14816
rect 1104 14714 38272 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38272 14714
rect 1104 14640 38272 14662
rect 3145 14603 3203 14609
rect 3145 14569 3157 14603
rect 3191 14600 3203 14603
rect 3234 14600 3240 14612
rect 3191 14572 3240 14600
rect 3191 14569 3203 14572
rect 3145 14563 3203 14569
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 3602 14560 3608 14612
rect 3660 14560 3666 14612
rect 4062 14560 4068 14612
rect 4120 14560 4126 14612
rect 7377 14603 7435 14609
rect 7377 14569 7389 14603
rect 7423 14600 7435 14603
rect 7466 14600 7472 14612
rect 7423 14572 7472 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 7466 14560 7472 14572
rect 7524 14560 7530 14612
rect 13449 14603 13507 14609
rect 13449 14569 13461 14603
rect 13495 14600 13507 14603
rect 14090 14600 14096 14612
rect 13495 14572 14096 14600
rect 13495 14569 13507 14572
rect 13449 14563 13507 14569
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 15838 14560 15844 14612
rect 15896 14600 15902 14612
rect 16577 14603 16635 14609
rect 16577 14600 16589 14603
rect 15896 14572 16589 14600
rect 15896 14560 15902 14572
rect 16577 14569 16589 14572
rect 16623 14569 16635 14603
rect 16577 14563 16635 14569
rect 17034 14560 17040 14612
rect 17092 14560 17098 14612
rect 17402 14560 17408 14612
rect 17460 14600 17466 14612
rect 19613 14603 19671 14609
rect 19613 14600 19625 14603
rect 17460 14572 19625 14600
rect 17460 14560 17466 14572
rect 19613 14569 19625 14572
rect 19659 14569 19671 14603
rect 19613 14563 19671 14569
rect 22278 14560 22284 14612
rect 22336 14560 22342 14612
rect 23106 14560 23112 14612
rect 23164 14600 23170 14612
rect 23753 14603 23811 14609
rect 23753 14600 23765 14603
rect 23164 14572 23765 14600
rect 23164 14560 23170 14572
rect 23753 14569 23765 14572
rect 23799 14600 23811 14603
rect 26418 14600 26424 14612
rect 23799 14572 26424 14600
rect 23799 14569 23811 14572
rect 23753 14563 23811 14569
rect 26418 14560 26424 14572
rect 26476 14560 26482 14612
rect 28350 14560 28356 14612
rect 28408 14600 28414 14612
rect 31941 14603 31999 14609
rect 28408 14572 31800 14600
rect 28408 14560 28414 14572
rect 1394 14356 1400 14408
rect 1452 14356 1458 14408
rect 3620 14396 3648 14560
rect 13814 14492 13820 14544
rect 13872 14532 13878 14544
rect 13872 14504 17356 14532
rect 13872 14492 13878 14504
rect 3694 14424 3700 14476
rect 3752 14464 3758 14476
rect 3752 14436 7144 14464
rect 3752 14424 3758 14436
rect 4065 14399 4123 14405
rect 4065 14396 4077 14399
rect 3620 14368 4077 14396
rect 4065 14365 4077 14368
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14396 4307 14399
rect 4614 14396 4620 14408
rect 4295 14368 4620 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 5626 14356 5632 14408
rect 5684 14356 5690 14408
rect 7116 14396 7144 14436
rect 8570 14424 8576 14476
rect 8628 14464 8634 14476
rect 10137 14467 10195 14473
rect 8628 14436 9352 14464
rect 8628 14424 8634 14436
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 7116 14368 8953 14396
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 8941 14359 8999 14365
rect 9030 14356 9036 14408
rect 9088 14396 9094 14408
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 9088 14368 9137 14396
rect 9088 14356 9094 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9214 14356 9220 14408
rect 9272 14356 9278 14408
rect 9324 14405 9352 14436
rect 10137 14433 10149 14467
rect 10183 14464 10195 14467
rect 10226 14464 10232 14476
rect 10183 14436 10232 14464
rect 10183 14433 10195 14436
rect 10137 14427 10195 14433
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 11885 14467 11943 14473
rect 11885 14433 11897 14467
rect 11931 14464 11943 14467
rect 12158 14464 12164 14476
rect 11931 14436 12164 14464
rect 11931 14433 11943 14436
rect 11885 14427 11943 14433
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 12618 14424 12624 14476
rect 12676 14464 12682 14476
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 12676 14436 12817 14464
rect 12676 14424 12682 14436
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 12989 14467 13047 14473
rect 12989 14433 13001 14467
rect 13035 14464 13047 14467
rect 14366 14464 14372 14476
rect 13035 14436 14372 14464
rect 13035 14433 13047 14436
rect 12989 14427 13047 14433
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 15010 14424 15016 14476
rect 15068 14464 15074 14476
rect 15565 14467 15623 14473
rect 15565 14464 15577 14467
rect 15068 14436 15577 14464
rect 15068 14424 15074 14436
rect 15565 14433 15577 14436
rect 15611 14433 15623 14467
rect 17328 14464 17356 14504
rect 17770 14492 17776 14544
rect 17828 14532 17834 14544
rect 20162 14532 20168 14544
rect 17828 14504 20168 14532
rect 17828 14492 17834 14504
rect 15565 14427 15623 14433
rect 16408 14436 17080 14464
rect 17328 14436 17632 14464
rect 9309 14399 9367 14405
rect 9309 14365 9321 14399
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 9858 14356 9864 14408
rect 9916 14356 9922 14408
rect 12406 14368 13124 14396
rect 1670 14288 1676 14340
rect 1728 14288 1734 14340
rect 2958 14328 2964 14340
rect 2898 14300 2964 14328
rect 2958 14288 2964 14300
rect 3016 14288 3022 14340
rect 5902 14288 5908 14340
rect 5960 14288 5966 14340
rect 6914 14288 6920 14340
rect 6972 14288 6978 14340
rect 9582 14288 9588 14340
rect 9640 14288 9646 14340
rect 12250 14328 12256 14340
rect 11362 14300 12256 14328
rect 12250 14288 12256 14300
rect 12308 14288 12314 14340
rect 8662 14220 8668 14272
rect 8720 14260 8726 14272
rect 12406 14260 12434 14368
rect 13096 14269 13124 14368
rect 15286 14356 15292 14408
rect 15344 14356 15350 14408
rect 15580 14328 15608 14427
rect 16408 14408 16436 14436
rect 16390 14356 16396 14408
rect 16448 14356 16454 14408
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14396 16635 14399
rect 16666 14396 16672 14408
rect 16623 14368 16672 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 16758 14356 16764 14408
rect 16816 14356 16822 14408
rect 17052 14405 17080 14436
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14365 17095 14399
rect 17215 14399 17273 14405
rect 17215 14396 17227 14399
rect 17037 14359 17095 14365
rect 17144 14368 17227 14396
rect 16942 14328 16948 14340
rect 15580 14300 16948 14328
rect 16942 14288 16948 14300
rect 17000 14288 17006 14340
rect 8720 14232 12434 14260
rect 13081 14263 13139 14269
rect 8720 14220 8726 14232
rect 13081 14229 13093 14263
rect 13127 14260 13139 14263
rect 13998 14260 14004 14272
rect 13127 14232 14004 14260
rect 13127 14229 13139 14232
rect 13081 14223 13139 14229
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 14274 14220 14280 14272
rect 14332 14260 14338 14272
rect 15746 14260 15752 14272
rect 14332 14232 15752 14260
rect 14332 14220 14338 14232
rect 15746 14220 15752 14232
rect 15804 14220 15810 14272
rect 15930 14220 15936 14272
rect 15988 14260 15994 14272
rect 17144 14260 17172 14368
rect 17215 14365 17227 14368
rect 17261 14365 17273 14399
rect 17215 14359 17273 14365
rect 17313 14399 17371 14405
rect 17313 14365 17325 14399
rect 17359 14396 17371 14399
rect 17604 14396 17632 14436
rect 17678 14424 17684 14476
rect 17736 14464 17742 14476
rect 18049 14467 18107 14473
rect 18049 14464 18061 14467
rect 17736 14436 18061 14464
rect 17736 14424 17742 14436
rect 18049 14433 18061 14436
rect 18095 14433 18107 14467
rect 18049 14427 18107 14433
rect 17957 14399 18015 14405
rect 17957 14396 17969 14399
rect 17359 14368 17448 14396
rect 17604 14368 17969 14396
rect 17359 14365 17371 14368
rect 17313 14359 17371 14365
rect 17420 14340 17448 14368
rect 17957 14365 17969 14368
rect 18003 14365 18015 14399
rect 17957 14359 18015 14365
rect 17402 14288 17408 14340
rect 17460 14288 17466 14340
rect 18064 14328 18092 14427
rect 18156 14405 18184 14504
rect 20162 14492 20168 14504
rect 20220 14492 20226 14544
rect 20530 14492 20536 14544
rect 20588 14492 20594 14544
rect 20622 14492 20628 14544
rect 20680 14532 20686 14544
rect 20680 14504 21312 14532
rect 20680 14492 20686 14504
rect 20548 14464 20576 14492
rect 20993 14467 21051 14473
rect 20993 14464 21005 14467
rect 20548 14436 21005 14464
rect 20993 14433 21005 14436
rect 21039 14433 21051 14467
rect 20993 14427 21051 14433
rect 18141 14399 18199 14405
rect 18141 14365 18153 14399
rect 18187 14365 18199 14399
rect 18141 14359 18199 14365
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14365 19947 14399
rect 19889 14359 19947 14365
rect 19245 14331 19303 14337
rect 19245 14328 19257 14331
rect 18064 14300 19257 14328
rect 19245 14297 19257 14300
rect 19291 14297 19303 14331
rect 19904 14328 19932 14359
rect 20070 14356 20076 14408
rect 20128 14396 20134 14408
rect 20257 14399 20315 14405
rect 20257 14396 20269 14399
rect 20128 14368 20269 14396
rect 20128 14356 20134 14368
rect 20257 14365 20269 14368
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 20533 14399 20591 14405
rect 20533 14365 20545 14399
rect 20579 14365 20591 14399
rect 20533 14359 20591 14365
rect 20438 14328 20444 14340
rect 19904 14300 20444 14328
rect 19245 14291 19303 14297
rect 20438 14288 20444 14300
rect 20496 14328 20502 14340
rect 20548 14328 20576 14359
rect 21082 14356 21088 14408
rect 21140 14356 21146 14408
rect 21284 14405 21312 14504
rect 22738 14492 22744 14544
rect 22796 14532 22802 14544
rect 29178 14532 29184 14544
rect 22796 14504 29184 14532
rect 22796 14492 22802 14504
rect 29178 14492 29184 14504
rect 29236 14492 29242 14544
rect 31018 14492 31024 14544
rect 31076 14492 31082 14544
rect 31570 14532 31576 14544
rect 31404 14504 31576 14532
rect 21637 14467 21695 14473
rect 21637 14433 21649 14467
rect 21683 14464 21695 14467
rect 22094 14464 22100 14476
rect 21683 14436 22100 14464
rect 21683 14433 21695 14436
rect 21637 14427 21695 14433
rect 22094 14424 22100 14436
rect 22152 14464 22158 14476
rect 22278 14464 22284 14476
rect 22152 14436 22284 14464
rect 22152 14424 22158 14436
rect 22278 14424 22284 14436
rect 22336 14464 22342 14476
rect 22336 14436 22692 14464
rect 22336 14424 22342 14436
rect 22664 14405 22692 14436
rect 23198 14424 23204 14476
rect 23256 14464 23262 14476
rect 23293 14467 23351 14473
rect 23293 14464 23305 14467
rect 23256 14436 23305 14464
rect 23256 14424 23262 14436
rect 23293 14433 23305 14436
rect 23339 14433 23351 14467
rect 23293 14427 23351 14433
rect 23385 14467 23443 14473
rect 23385 14433 23397 14467
rect 23431 14464 23443 14467
rect 30193 14467 30251 14473
rect 23431 14436 24164 14464
rect 23431 14433 23443 14436
rect 23385 14427 23443 14433
rect 21269 14399 21327 14405
rect 21269 14365 21281 14399
rect 21315 14365 21327 14399
rect 21269 14359 21327 14365
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14365 22063 14399
rect 22005 14359 22063 14365
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14365 22707 14399
rect 22649 14359 22707 14365
rect 20496 14300 20576 14328
rect 21100 14328 21128 14356
rect 21818 14328 21824 14340
rect 21100 14300 21824 14328
rect 20496 14288 20502 14300
rect 21818 14288 21824 14300
rect 21876 14328 21882 14340
rect 22020 14328 22048 14359
rect 22830 14356 22836 14408
rect 22888 14356 22894 14408
rect 23308 14396 23336 14427
rect 24136 14408 24164 14436
rect 30193 14433 30205 14467
rect 30239 14464 30251 14467
rect 30650 14464 30656 14476
rect 30239 14436 30656 14464
rect 30239 14433 30251 14436
rect 30193 14427 30251 14433
rect 30650 14424 30656 14436
rect 30708 14424 30714 14476
rect 30834 14424 30840 14476
rect 30892 14424 30898 14476
rect 23474 14396 23480 14408
rect 23308 14368 23480 14396
rect 23474 14356 23480 14368
rect 23532 14356 23538 14408
rect 23569 14399 23627 14405
rect 23569 14365 23581 14399
rect 23615 14365 23627 14399
rect 23569 14359 23627 14365
rect 21876 14300 22048 14328
rect 22848 14328 22876 14356
rect 23198 14328 23204 14340
rect 22848 14300 23204 14328
rect 21876 14288 21882 14300
rect 23198 14288 23204 14300
rect 23256 14328 23262 14340
rect 23584 14328 23612 14359
rect 24118 14356 24124 14408
rect 24176 14356 24182 14408
rect 25498 14356 25504 14408
rect 25556 14396 25562 14408
rect 27154 14396 27160 14408
rect 25556 14368 27160 14396
rect 25556 14356 25562 14368
rect 27154 14356 27160 14368
rect 27212 14356 27218 14408
rect 30377 14399 30435 14405
rect 30377 14365 30389 14399
rect 30423 14396 30435 14399
rect 30852 14396 30880 14424
rect 31036 14396 31064 14492
rect 31404 14405 31432 14504
rect 31570 14492 31576 14504
rect 31628 14492 31634 14544
rect 31662 14464 31668 14476
rect 31496 14436 31668 14464
rect 31496 14405 31524 14436
rect 31662 14424 31668 14436
rect 31720 14424 31726 14476
rect 31772 14405 31800 14572
rect 31941 14569 31953 14603
rect 31987 14600 31999 14603
rect 32950 14600 32956 14612
rect 31987 14572 32956 14600
rect 31987 14569 31999 14572
rect 31941 14563 31999 14569
rect 32950 14560 32956 14572
rect 33008 14560 33014 14612
rect 31205 14399 31263 14405
rect 31205 14396 31217 14399
rect 30423 14368 30972 14396
rect 31036 14368 31217 14396
rect 30423 14365 30435 14368
rect 30377 14359 30435 14365
rect 23256 14300 23612 14328
rect 30561 14331 30619 14337
rect 23256 14288 23262 14300
rect 30561 14297 30573 14331
rect 30607 14328 30619 14331
rect 30653 14331 30711 14337
rect 30653 14328 30665 14331
rect 30607 14300 30665 14328
rect 30607 14297 30619 14300
rect 30561 14291 30619 14297
rect 30653 14297 30665 14300
rect 30699 14297 30711 14331
rect 30653 14291 30711 14297
rect 30742 14288 30748 14340
rect 30800 14328 30806 14340
rect 30837 14331 30895 14337
rect 30837 14328 30849 14331
rect 30800 14300 30849 14328
rect 30800 14288 30806 14300
rect 30837 14297 30849 14300
rect 30883 14297 30895 14331
rect 30944 14328 30972 14368
rect 31205 14365 31217 14368
rect 31251 14365 31263 14399
rect 31205 14359 31263 14365
rect 31389 14399 31447 14405
rect 31389 14365 31401 14399
rect 31435 14365 31447 14399
rect 31389 14359 31447 14365
rect 31481 14399 31539 14405
rect 31481 14365 31493 14399
rect 31527 14365 31539 14399
rect 31481 14359 31539 14365
rect 31573 14399 31631 14405
rect 31573 14365 31585 14399
rect 31619 14396 31631 14399
rect 31757 14399 31815 14405
rect 31619 14368 31708 14396
rect 31619 14365 31631 14368
rect 31573 14359 31631 14365
rect 30944 14300 31248 14328
rect 30837 14291 30895 14297
rect 31220 14272 31248 14300
rect 19334 14260 19340 14272
rect 15988 14232 19340 14260
rect 15988 14220 15994 14232
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 19622 14263 19680 14269
rect 19622 14229 19634 14263
rect 19668 14260 19680 14263
rect 19978 14260 19984 14272
rect 19668 14232 19984 14260
rect 19668 14229 19680 14232
rect 19622 14223 19680 14229
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 22830 14220 22836 14272
rect 22888 14260 22894 14272
rect 25130 14260 25136 14272
rect 22888 14232 25136 14260
rect 22888 14220 22894 14232
rect 25130 14220 25136 14232
rect 25188 14220 25194 14272
rect 25774 14220 25780 14272
rect 25832 14260 25838 14272
rect 26234 14260 26240 14272
rect 25832 14232 26240 14260
rect 25832 14220 25838 14232
rect 26234 14220 26240 14232
rect 26292 14260 26298 14272
rect 27062 14260 27068 14272
rect 26292 14232 27068 14260
rect 26292 14220 26298 14232
rect 27062 14220 27068 14232
rect 27120 14220 27126 14272
rect 29270 14220 29276 14272
rect 29328 14260 29334 14272
rect 30190 14260 30196 14272
rect 29328 14232 30196 14260
rect 29328 14220 29334 14232
rect 30190 14220 30196 14232
rect 30248 14220 30254 14272
rect 30374 14220 30380 14272
rect 30432 14260 30438 14272
rect 31021 14263 31079 14269
rect 31021 14260 31033 14263
rect 30432 14232 31033 14260
rect 30432 14220 30438 14232
rect 31021 14229 31033 14232
rect 31067 14229 31079 14263
rect 31021 14223 31079 14229
rect 31202 14220 31208 14272
rect 31260 14220 31266 14272
rect 31386 14220 31392 14272
rect 31444 14260 31450 14272
rect 31680 14260 31708 14368
rect 31757 14365 31769 14399
rect 31803 14365 31815 14399
rect 31757 14359 31815 14365
rect 33778 14260 33784 14272
rect 31444 14232 33784 14260
rect 31444 14220 31450 14232
rect 33778 14220 33784 14232
rect 33836 14260 33842 14272
rect 34054 14260 34060 14272
rect 33836 14232 34060 14260
rect 33836 14220 33842 14232
rect 34054 14220 34060 14232
rect 34112 14220 34118 14272
rect 1104 14170 38272 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38272 14170
rect 1104 14096 38272 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 1949 14059 2007 14065
rect 1949 14056 1961 14059
rect 1728 14028 1961 14056
rect 1728 14016 1734 14028
rect 1949 14025 1961 14028
rect 1995 14025 2007 14059
rect 1949 14019 2007 14025
rect 2498 14016 2504 14068
rect 2556 14016 2562 14068
rect 5902 14016 5908 14068
rect 5960 14056 5966 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 5960 14028 6377 14056
rect 5960 14016 5966 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 6365 14019 6423 14025
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14025 6699 14059
rect 6641 14019 6699 14025
rect 7009 14059 7067 14065
rect 7009 14025 7021 14059
rect 7055 14056 7067 14059
rect 8662 14056 8668 14068
rect 7055 14028 8668 14056
rect 7055 14025 7067 14028
rect 7009 14019 7067 14025
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 2516 13920 2544 14016
rect 2179 13892 2544 13920
rect 6549 13923 6607 13929
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 6549 13889 6561 13923
rect 6595 13920 6607 13923
rect 6656 13920 6684 14019
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 13814 14056 13820 14068
rect 12032 14028 13820 14056
rect 12032 14016 12038 14028
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 16942 14016 16948 14068
rect 17000 14056 17006 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17000 14028 17785 14056
rect 17000 14016 17006 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 17773 14019 17831 14025
rect 17865 14059 17923 14065
rect 17865 14025 17877 14059
rect 17911 14056 17923 14059
rect 19426 14056 19432 14068
rect 17911 14028 19432 14056
rect 17911 14025 17923 14028
rect 17865 14019 17923 14025
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 19797 14059 19855 14065
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 21082 14056 21088 14068
rect 19843 14028 21088 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 21266 14016 21272 14068
rect 21324 14016 21330 14068
rect 22186 14016 22192 14068
rect 22244 14056 22250 14068
rect 22830 14056 22836 14068
rect 22244 14028 22836 14056
rect 22244 14016 22250 14028
rect 22830 14016 22836 14028
rect 22888 14016 22894 14068
rect 23477 14059 23535 14065
rect 23477 14025 23489 14059
rect 23523 14056 23535 14059
rect 23523 14028 25912 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 7101 13991 7159 13997
rect 7101 13957 7113 13991
rect 7147 13988 7159 13991
rect 7466 13988 7472 14000
rect 7147 13960 7472 13988
rect 7147 13957 7159 13960
rect 7101 13951 7159 13957
rect 7466 13948 7472 13960
rect 7524 13948 7530 14000
rect 8294 13948 8300 14000
rect 8352 13988 8358 14000
rect 10134 13988 10140 14000
rect 8352 13960 10140 13988
rect 8352 13948 8358 13960
rect 6595 13892 6684 13920
rect 6595 13889 6607 13892
rect 6549 13883 6607 13889
rect 1486 13812 1492 13864
rect 1544 13812 1550 13864
rect 1780 13852 1808 13883
rect 8386 13880 8392 13932
rect 8444 13880 8450 13932
rect 8496 13929 8524 13960
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 17221 13991 17279 13997
rect 14660 13960 16804 13988
rect 14660 13932 14688 13960
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 9950 13880 9956 13932
rect 10008 13920 10014 13932
rect 12802 13920 12808 13932
rect 10008 13892 12808 13920
rect 10008 13880 10014 13892
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 13354 13880 13360 13932
rect 13412 13880 13418 13932
rect 14642 13880 14648 13932
rect 14700 13880 14706 13932
rect 15194 13880 15200 13932
rect 15252 13920 15258 13932
rect 16776 13929 16804 13960
rect 17221 13957 17233 13991
rect 17267 13988 17279 13991
rect 17310 13988 17316 14000
rect 17267 13960 17316 13988
rect 17267 13957 17279 13960
rect 17221 13951 17279 13957
rect 17310 13948 17316 13960
rect 17368 13948 17374 14000
rect 20070 13988 20076 14000
rect 19628 13960 20076 13988
rect 19628 13932 19656 13960
rect 20070 13948 20076 13960
rect 20128 13988 20134 14000
rect 20128 13960 20392 13988
rect 20128 13948 20134 13960
rect 15289 13923 15347 13929
rect 15289 13920 15301 13923
rect 15252 13892 15301 13920
rect 15252 13880 15258 13892
rect 15289 13889 15301 13892
rect 15335 13920 15347 13923
rect 16209 13923 16267 13929
rect 16209 13920 16221 13923
rect 15335 13892 16221 13920
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 16209 13889 16221 13892
rect 16255 13920 16267 13923
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16255 13892 16681 13920
rect 16255 13889 16267 13892
rect 16209 13883 16267 13889
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 16761 13923 16819 13929
rect 16761 13889 16773 13923
rect 16807 13920 16819 13923
rect 17126 13920 17132 13932
rect 16807 13892 17132 13920
rect 16807 13889 16819 13892
rect 16761 13883 16819 13889
rect 17126 13880 17132 13892
rect 17184 13920 17190 13932
rect 17402 13920 17408 13932
rect 17184 13892 17408 13920
rect 17184 13880 17190 13892
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 19610 13920 19616 13932
rect 17880 13892 19616 13920
rect 5534 13852 5540 13864
rect 1780 13824 5540 13852
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 7190 13812 7196 13864
rect 7248 13812 7254 13864
rect 13372 13852 13400 13880
rect 15565 13855 15623 13861
rect 15565 13852 15577 13855
rect 13372 13824 15577 13852
rect 15565 13821 15577 13824
rect 15611 13852 15623 13855
rect 16850 13852 16856 13864
rect 15611 13824 16856 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 16850 13812 16856 13824
rect 16908 13852 16914 13864
rect 17880 13852 17908 13892
rect 19610 13880 19616 13892
rect 19668 13880 19674 13932
rect 19702 13880 19708 13932
rect 19760 13880 19766 13932
rect 20257 13923 20315 13929
rect 20257 13920 20269 13923
rect 19812 13892 20269 13920
rect 16908 13824 17908 13852
rect 17957 13855 18015 13861
rect 16908 13812 16914 13824
rect 17957 13821 17969 13855
rect 18003 13821 18015 13855
rect 17957 13815 18015 13821
rect 10962 13744 10968 13796
rect 11020 13784 11026 13796
rect 17972 13784 18000 13815
rect 11020 13756 18000 13784
rect 11020 13744 11026 13756
rect 18414 13744 18420 13796
rect 18472 13784 18478 13796
rect 19150 13784 19156 13796
rect 18472 13756 19156 13784
rect 18472 13744 18478 13756
rect 19150 13744 19156 13756
rect 19208 13744 19214 13796
rect 9398 13676 9404 13728
rect 9456 13716 9462 13728
rect 12526 13716 12532 13728
rect 9456 13688 12532 13716
rect 9456 13676 9462 13688
rect 12526 13676 12532 13688
rect 12584 13676 12590 13728
rect 15013 13719 15071 13725
rect 15013 13685 15025 13719
rect 15059 13716 15071 13719
rect 15562 13716 15568 13728
rect 15059 13688 15568 13716
rect 15059 13685 15071 13688
rect 15013 13679 15071 13685
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 17402 13676 17408 13728
rect 17460 13676 17466 13728
rect 17862 13676 17868 13728
rect 17920 13716 17926 13728
rect 19426 13716 19432 13728
rect 17920 13688 19432 13716
rect 17920 13676 17926 13688
rect 19426 13676 19432 13688
rect 19484 13716 19490 13728
rect 19812 13716 19840 13892
rect 20257 13889 20269 13892
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 20364 13784 20392 13960
rect 20530 13948 20536 14000
rect 20588 13988 20594 14000
rect 20588 13960 21128 13988
rect 20588 13948 20594 13960
rect 20438 13880 20444 13932
rect 20496 13920 20502 13932
rect 20625 13923 20683 13929
rect 20625 13920 20637 13923
rect 20496 13892 20637 13920
rect 20496 13880 20502 13892
rect 20625 13889 20637 13892
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 20640 13852 20668 13883
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 21100 13929 21128 13960
rect 20901 13923 20959 13929
rect 20901 13920 20913 13923
rect 20772 13892 20913 13920
rect 20772 13880 20778 13892
rect 20901 13889 20913 13892
rect 20947 13889 20959 13923
rect 20901 13883 20959 13889
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13889 21235 13923
rect 21284 13919 21312 14016
rect 23198 13948 23204 14000
rect 23256 13988 23262 14000
rect 25409 13991 25467 13997
rect 25409 13988 25421 13991
rect 23256 13960 24440 13988
rect 23256 13948 23262 13960
rect 21177 13883 21235 13889
rect 21270 13913 21328 13919
rect 21192 13852 21220 13883
rect 21270 13879 21282 13913
rect 21316 13879 21328 13913
rect 21818 13880 21824 13932
rect 21876 13920 21882 13932
rect 22097 13923 22155 13929
rect 22097 13920 22109 13923
rect 21876 13892 22109 13920
rect 21876 13880 21882 13892
rect 22097 13889 22109 13892
rect 22143 13889 22155 13923
rect 22097 13883 22155 13889
rect 22281 13923 22339 13929
rect 22281 13889 22293 13923
rect 22327 13920 22339 13923
rect 22649 13923 22707 13929
rect 22649 13920 22661 13923
rect 22327 13892 22661 13920
rect 22327 13889 22339 13892
rect 22281 13883 22339 13889
rect 22649 13889 22661 13892
rect 22695 13920 22707 13923
rect 24118 13920 24124 13932
rect 22695 13892 24124 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 24118 13880 24124 13892
rect 24176 13880 24182 13932
rect 24412 13929 24440 13960
rect 24872 13960 25421 13988
rect 24397 13923 24455 13929
rect 24397 13889 24409 13923
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 24762 13880 24768 13932
rect 24820 13880 24826 13932
rect 24872 13929 24900 13960
rect 25409 13957 25421 13960
rect 25455 13957 25467 13991
rect 25774 13988 25780 14000
rect 25409 13951 25467 13957
rect 25700 13960 25780 13988
rect 24857 13923 24915 13929
rect 24857 13889 24869 13923
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 25038 13880 25044 13932
rect 25096 13880 25102 13932
rect 25130 13880 25136 13932
rect 25188 13880 25194 13932
rect 25700 13929 25728 13960
rect 25774 13948 25780 13960
rect 25832 13948 25838 14000
rect 25884 13929 25912 14028
rect 26326 14016 26332 14068
rect 26384 14056 26390 14068
rect 26384 14028 26556 14056
rect 26384 14016 26390 14028
rect 26421 13991 26479 13997
rect 26421 13988 26433 13991
rect 25976 13960 26433 13988
rect 25976 13929 26004 13960
rect 26421 13957 26433 13960
rect 26467 13957 26479 13991
rect 26421 13951 26479 13957
rect 25593 13923 25651 13929
rect 25593 13889 25605 13923
rect 25639 13889 25651 13923
rect 25593 13883 25651 13889
rect 25685 13923 25743 13929
rect 25685 13889 25697 13923
rect 25731 13889 25743 13923
rect 25685 13883 25743 13889
rect 25869 13923 25927 13929
rect 25869 13889 25881 13923
rect 25915 13889 25927 13923
rect 25869 13883 25927 13889
rect 25961 13923 26019 13929
rect 25961 13889 25973 13923
rect 26007 13889 26019 13923
rect 25961 13883 26019 13889
rect 26053 13923 26111 13929
rect 26053 13889 26065 13923
rect 26099 13889 26111 13923
rect 26053 13883 26111 13889
rect 21270 13873 21328 13879
rect 20640 13824 21220 13852
rect 21284 13784 21312 13873
rect 21913 13855 21971 13861
rect 21913 13821 21925 13855
rect 21959 13821 21971 13855
rect 21913 13815 21971 13821
rect 20364 13756 21312 13784
rect 21358 13744 21364 13796
rect 21416 13784 21422 13796
rect 21545 13787 21603 13793
rect 21545 13784 21557 13787
rect 21416 13756 21557 13784
rect 21416 13744 21422 13756
rect 21545 13753 21557 13756
rect 21591 13784 21603 13787
rect 21928 13784 21956 13815
rect 22370 13812 22376 13864
rect 22428 13852 22434 13864
rect 22465 13855 22523 13861
rect 22465 13852 22477 13855
rect 22428 13824 22477 13852
rect 22428 13812 22434 13824
rect 22465 13821 22477 13824
rect 22511 13821 22523 13855
rect 22465 13815 22523 13821
rect 21591 13756 21956 13784
rect 21591 13753 21603 13756
rect 21545 13747 21603 13753
rect 19484 13688 19840 13716
rect 22480 13716 22508 13815
rect 22554 13812 22560 13864
rect 22612 13812 22618 13864
rect 22738 13812 22744 13864
rect 22796 13852 22802 13864
rect 23017 13855 23075 13861
rect 23017 13852 23029 13855
rect 22796 13824 23029 13852
rect 22796 13812 22802 13824
rect 23017 13821 23029 13824
rect 23063 13821 23075 13855
rect 23017 13815 23075 13821
rect 23109 13855 23167 13861
rect 23109 13821 23121 13855
rect 23155 13821 23167 13855
rect 23109 13815 23167 13821
rect 22572 13784 22600 13812
rect 22922 13784 22928 13796
rect 22572 13756 22928 13784
rect 22922 13744 22928 13756
rect 22980 13784 22986 13796
rect 23124 13784 23152 13815
rect 23198 13812 23204 13864
rect 23256 13812 23262 13864
rect 23293 13855 23351 13861
rect 23293 13821 23305 13855
rect 23339 13821 23351 13855
rect 23293 13815 23351 13821
rect 22980 13756 23152 13784
rect 22980 13744 22986 13756
rect 22554 13716 22560 13728
rect 22480 13688 22560 13716
rect 19484 13676 19490 13688
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 22738 13676 22744 13728
rect 22796 13716 22802 13728
rect 23308 13716 23336 13815
rect 23474 13812 23480 13864
rect 23532 13852 23538 13864
rect 23658 13852 23664 13864
rect 23532 13824 23664 13852
rect 23532 13812 23538 13824
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 23842 13812 23848 13864
rect 23900 13852 23906 13864
rect 25608 13852 25636 13883
rect 26068 13852 26096 13883
rect 26142 13880 26148 13932
rect 26200 13920 26206 13932
rect 26528 13929 26556 14028
rect 27246 14016 27252 14068
rect 27304 14016 27310 14068
rect 28442 14016 28448 14068
rect 28500 14056 28506 14068
rect 29089 14059 29147 14065
rect 29089 14056 29101 14059
rect 28500 14028 29101 14056
rect 28500 14016 28506 14028
rect 29089 14025 29101 14028
rect 29135 14025 29147 14059
rect 29089 14019 29147 14025
rect 29178 14016 29184 14068
rect 29236 14056 29242 14068
rect 30834 14056 30840 14068
rect 29236 14028 30840 14056
rect 29236 14016 29242 14028
rect 30834 14016 30840 14028
rect 30892 14016 30898 14068
rect 31389 14059 31447 14065
rect 31389 14025 31401 14059
rect 31435 14056 31447 14059
rect 31478 14056 31484 14068
rect 31435 14028 31484 14056
rect 31435 14025 31447 14028
rect 31389 14019 31447 14025
rect 31478 14016 31484 14028
rect 31536 14016 31542 14068
rect 32858 14016 32864 14068
rect 32916 14016 32922 14068
rect 27264 13988 27292 14016
rect 26804 13960 27292 13988
rect 26804 13929 26832 13960
rect 26237 13923 26295 13929
rect 26237 13920 26249 13923
rect 26200 13892 26249 13920
rect 26200 13880 26206 13892
rect 26237 13889 26249 13892
rect 26283 13889 26295 13923
rect 26237 13883 26295 13889
rect 26329 13923 26387 13929
rect 26329 13889 26341 13923
rect 26375 13889 26387 13923
rect 26329 13883 26387 13889
rect 26513 13923 26571 13929
rect 26513 13889 26525 13923
rect 26559 13889 26571 13923
rect 26513 13883 26571 13889
rect 26605 13923 26663 13929
rect 26605 13889 26617 13923
rect 26651 13889 26663 13923
rect 26605 13883 26663 13889
rect 26789 13923 26847 13929
rect 26789 13889 26801 13923
rect 26835 13889 26847 13923
rect 26789 13883 26847 13889
rect 26344 13852 26372 13883
rect 23900 13824 25636 13852
rect 25700 13824 26096 13852
rect 26252 13824 26372 13852
rect 26620 13852 26648 13883
rect 27062 13880 27068 13932
rect 27120 13880 27126 13932
rect 27264 13929 27292 13960
rect 27798 13948 27804 14000
rect 27856 13988 27862 14000
rect 32876 13988 32904 14016
rect 27856 13960 30236 13988
rect 27856 13948 27862 13960
rect 27249 13923 27307 13929
rect 27249 13889 27261 13923
rect 27295 13889 27307 13923
rect 27249 13883 27307 13889
rect 28074 13880 28080 13932
rect 28132 13920 28138 13932
rect 28810 13920 28816 13932
rect 28132 13892 28816 13920
rect 28132 13880 28138 13892
rect 28810 13880 28816 13892
rect 28868 13880 28874 13932
rect 29089 13923 29147 13929
rect 29089 13889 29101 13923
rect 29135 13889 29147 13923
rect 29089 13883 29147 13889
rect 27080 13852 27108 13880
rect 26620 13824 27108 13852
rect 28905 13855 28963 13861
rect 23900 13812 23906 13824
rect 24394 13744 24400 13796
rect 24452 13744 24458 13796
rect 25317 13787 25375 13793
rect 25317 13753 25329 13787
rect 25363 13784 25375 13787
rect 25498 13784 25504 13796
rect 25363 13756 25504 13784
rect 25363 13753 25375 13756
rect 25317 13747 25375 13753
rect 25498 13744 25504 13756
rect 25556 13744 25562 13796
rect 24210 13716 24216 13728
rect 22796 13688 24216 13716
rect 22796 13676 22802 13688
rect 24210 13676 24216 13688
rect 24268 13716 24274 13728
rect 25700 13716 25728 13824
rect 26252 13784 26280 13824
rect 28905 13821 28917 13855
rect 28951 13852 28963 13855
rect 28994 13852 29000 13864
rect 28951 13824 29000 13852
rect 28951 13821 28963 13824
rect 28905 13815 28963 13821
rect 28994 13812 29000 13824
rect 29052 13812 29058 13864
rect 27246 13784 27252 13796
rect 26252 13756 27252 13784
rect 26252 13728 26280 13756
rect 27246 13744 27252 13756
rect 27304 13744 27310 13796
rect 29104 13784 29132 13883
rect 29178 13880 29184 13932
rect 29236 13920 29242 13932
rect 30208 13929 30236 13960
rect 30300 13960 32812 13988
rect 32876 13960 33088 13988
rect 29273 13923 29331 13929
rect 29273 13920 29285 13923
rect 29236 13892 29285 13920
rect 29236 13880 29242 13892
rect 29273 13889 29285 13892
rect 29319 13889 29331 13923
rect 29273 13883 29331 13889
rect 30193 13923 30251 13929
rect 30193 13889 30205 13923
rect 30239 13889 30251 13923
rect 30193 13883 30251 13889
rect 30098 13852 30104 13864
rect 29288 13824 30104 13852
rect 29288 13796 29316 13824
rect 30098 13812 30104 13824
rect 30156 13852 30162 13864
rect 30300 13852 30328 13960
rect 30374 13880 30380 13932
rect 30432 13880 30438 13932
rect 30760 13929 30788 13960
rect 30745 13923 30803 13929
rect 30745 13889 30757 13923
rect 30791 13889 30803 13923
rect 30745 13883 30803 13889
rect 30834 13880 30840 13932
rect 30892 13880 30898 13932
rect 32784 13929 32812 13960
rect 30929 13923 30987 13929
rect 30929 13889 30941 13923
rect 30975 13920 30987 13923
rect 31941 13923 31999 13929
rect 31941 13920 31953 13923
rect 30975 13892 31953 13920
rect 30975 13889 30987 13892
rect 30929 13883 30987 13889
rect 31941 13889 31953 13892
rect 31987 13889 31999 13923
rect 31941 13883 31999 13889
rect 32769 13923 32827 13929
rect 32769 13889 32781 13923
rect 32815 13889 32827 13923
rect 32769 13883 32827 13889
rect 30156 13824 30328 13852
rect 30156 13812 30162 13824
rect 30466 13812 30472 13864
rect 30524 13812 30530 13864
rect 30561 13855 30619 13861
rect 30561 13821 30573 13855
rect 30607 13821 30619 13855
rect 30852 13852 30880 13880
rect 31665 13855 31723 13861
rect 30852 13824 31616 13852
rect 30561 13815 30619 13821
rect 28552 13756 29132 13784
rect 28552 13728 28580 13756
rect 24268 13688 25728 13716
rect 24268 13676 24274 13688
rect 25774 13676 25780 13728
rect 25832 13716 25838 13728
rect 26145 13719 26203 13725
rect 26145 13716 26157 13719
rect 25832 13688 26157 13716
rect 25832 13676 25838 13688
rect 26145 13685 26157 13688
rect 26191 13685 26203 13719
rect 26145 13679 26203 13685
rect 26234 13676 26240 13728
rect 26292 13676 26298 13728
rect 26694 13676 26700 13728
rect 26752 13716 26758 13728
rect 26789 13719 26847 13725
rect 26789 13716 26801 13719
rect 26752 13688 26801 13716
rect 26752 13676 26758 13688
rect 26789 13685 26801 13688
rect 26835 13685 26847 13719
rect 26789 13679 26847 13685
rect 27154 13676 27160 13728
rect 27212 13676 27218 13728
rect 28534 13676 28540 13728
rect 28592 13676 28598 13728
rect 29104 13716 29132 13756
rect 29270 13744 29276 13796
rect 29328 13744 29334 13796
rect 30576 13784 30604 13815
rect 30742 13784 30748 13796
rect 30576 13756 30748 13784
rect 30742 13744 30748 13756
rect 30800 13744 30806 13796
rect 31588 13784 31616 13824
rect 31665 13821 31677 13855
rect 31711 13852 31723 13855
rect 32398 13852 32404 13864
rect 31711 13824 32404 13852
rect 31711 13821 31723 13824
rect 31665 13815 31723 13821
rect 32398 13812 32404 13824
rect 32456 13812 32462 13864
rect 32784 13852 32812 13883
rect 32950 13880 32956 13932
rect 33008 13880 33014 13932
rect 33060 13929 33088 13960
rect 33045 13923 33103 13929
rect 33045 13889 33057 13923
rect 33091 13889 33103 13923
rect 33045 13883 33103 13889
rect 33226 13880 33232 13932
rect 33284 13880 33290 13932
rect 33502 13880 33508 13932
rect 33560 13880 33566 13932
rect 33520 13852 33548 13880
rect 32784 13824 33548 13852
rect 31588 13756 32628 13784
rect 32600 13728 32628 13756
rect 29454 13716 29460 13728
rect 29104 13688 29460 13716
rect 29454 13676 29460 13688
rect 29512 13676 29518 13728
rect 31846 13676 31852 13728
rect 31904 13676 31910 13728
rect 32582 13676 32588 13728
rect 32640 13676 32646 13728
rect 33134 13676 33140 13728
rect 33192 13716 33198 13728
rect 33229 13719 33287 13725
rect 33229 13716 33241 13719
rect 33192 13688 33241 13716
rect 33192 13676 33198 13688
rect 33229 13685 33241 13688
rect 33275 13685 33287 13719
rect 33229 13679 33287 13685
rect 1104 13626 38272 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38272 13626
rect 1104 13552 38272 13574
rect 4249 13515 4307 13521
rect 4249 13481 4261 13515
rect 4295 13512 4307 13515
rect 9030 13512 9036 13524
rect 4295 13484 9036 13512
rect 4295 13481 4307 13484
rect 4249 13475 4307 13481
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 10318 13472 10324 13524
rect 10376 13472 10382 13524
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 10468 13484 10517 13512
rect 10468 13472 10474 13484
rect 10505 13481 10517 13484
rect 10551 13481 10563 13515
rect 11238 13512 11244 13524
rect 10505 13475 10563 13481
rect 10612 13484 11244 13512
rect 9125 13447 9183 13453
rect 9125 13413 9137 13447
rect 9171 13413 9183 13447
rect 9125 13407 9183 13413
rect 1394 13336 1400 13388
rect 1452 13376 1458 13388
rect 4341 13379 4399 13385
rect 4341 13376 4353 13379
rect 1452 13348 4353 13376
rect 1452 13336 1458 13348
rect 4341 13345 4353 13348
rect 4387 13376 4399 13379
rect 5626 13376 5632 13388
rect 4387 13348 5632 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 5626 13336 5632 13348
rect 5684 13336 5690 13388
rect 6270 13336 6276 13388
rect 6328 13376 6334 13388
rect 6365 13379 6423 13385
rect 6365 13376 6377 13379
rect 6328 13348 6377 13376
rect 6328 13336 6334 13348
rect 6365 13345 6377 13348
rect 6411 13345 6423 13379
rect 6914 13376 6920 13388
rect 6365 13339 6423 13345
rect 6472 13348 6920 13376
rect 3326 13268 3332 13320
rect 3384 13308 3390 13320
rect 3786 13308 3792 13320
rect 3384 13280 3792 13308
rect 3384 13268 3390 13280
rect 3786 13268 3792 13280
rect 3844 13308 3850 13320
rect 3881 13311 3939 13317
rect 3881 13308 3893 13311
rect 3844 13280 3893 13308
rect 3844 13268 3850 13280
rect 3881 13277 3893 13280
rect 3927 13277 3939 13311
rect 3881 13271 3939 13277
rect 3970 13200 3976 13252
rect 4028 13240 4034 13252
rect 4065 13243 4123 13249
rect 4065 13240 4077 13243
rect 4028 13212 4077 13240
rect 4028 13200 4034 13212
rect 4065 13209 4077 13212
rect 4111 13209 4123 13243
rect 4065 13203 4123 13209
rect 4614 13200 4620 13252
rect 4672 13200 4678 13252
rect 5000 13212 5106 13240
rect 2958 13132 2964 13184
rect 3016 13172 3022 13184
rect 5000 13172 5028 13212
rect 6472 13172 6500 13348
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 7190 13336 7196 13388
rect 7248 13336 7254 13388
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13308 8815 13311
rect 9140 13308 9168 13407
rect 9582 13336 9588 13388
rect 9640 13336 9646 13388
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13376 9827 13379
rect 10336 13376 10364 13472
rect 9815 13348 10364 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 8803 13280 9168 13308
rect 8803 13277 8815 13280
rect 8757 13271 8815 13277
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 9600 13308 9628 13336
rect 9272 13280 10088 13308
rect 9272 13268 9278 13280
rect 6917 13243 6975 13249
rect 6917 13209 6929 13243
rect 6963 13240 6975 13243
rect 9950 13240 9956 13252
rect 6963 13212 9956 13240
rect 6963 13209 6975 13212
rect 6917 13203 6975 13209
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 10060 13240 10088 13280
rect 10134 13268 10140 13320
rect 10192 13268 10198 13320
rect 10612 13317 10640 13484
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 13814 13512 13820 13524
rect 12268 13484 13820 13512
rect 10965 13379 11023 13385
rect 10965 13345 10977 13379
rect 11011 13376 11023 13379
rect 11882 13376 11888 13388
rect 11011 13348 11888 13376
rect 11011 13345 11023 13348
rect 10965 13339 11023 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13277 10655 13311
rect 10597 13271 10655 13277
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 10244 13240 10272 13271
rect 10060 13212 10272 13240
rect 10704 13240 10732 13271
rect 12268 13252 12296 13484
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 14734 13472 14740 13524
rect 14792 13472 14798 13524
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 15381 13515 15439 13521
rect 15381 13512 15393 13515
rect 15344 13484 15393 13512
rect 15344 13472 15350 13484
rect 15381 13481 15393 13484
rect 15427 13481 15439 13515
rect 15381 13475 15439 13481
rect 16669 13515 16727 13521
rect 16669 13481 16681 13515
rect 16715 13512 16727 13515
rect 16758 13512 16764 13524
rect 16715 13484 16764 13512
rect 16715 13481 16727 13484
rect 16669 13475 16727 13481
rect 16758 13472 16764 13484
rect 16816 13512 16822 13524
rect 17218 13512 17224 13524
rect 16816 13484 17224 13512
rect 16816 13472 16822 13484
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 17862 13472 17868 13524
rect 17920 13472 17926 13524
rect 18414 13472 18420 13524
rect 18472 13472 18478 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 18524 13484 18889 13512
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 12897 13379 12955 13385
rect 12897 13376 12909 13379
rect 12676 13348 12909 13376
rect 12676 13336 12682 13348
rect 12897 13345 12909 13348
rect 12943 13345 12955 13379
rect 12897 13339 12955 13345
rect 13081 13379 13139 13385
rect 13081 13345 13093 13379
rect 13127 13376 13139 13379
rect 13354 13376 13360 13388
rect 13127 13348 13360 13376
rect 13127 13345 13139 13348
rect 13081 13339 13139 13345
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 14752 13376 14780 13472
rect 16850 13404 16856 13456
rect 16908 13404 16914 13456
rect 14752 13348 16804 13376
rect 12526 13268 12532 13320
rect 12584 13308 12590 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 12584 13280 13185 13308
rect 12584 13268 12590 13280
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 13817 13311 13875 13317
rect 13817 13308 13829 13311
rect 13173 13271 13231 13277
rect 13556 13280 13829 13308
rect 11146 13240 11152 13252
rect 10704 13212 11152 13240
rect 11146 13200 11152 13212
rect 11204 13200 11210 13252
rect 11241 13243 11299 13249
rect 11241 13209 11253 13243
rect 11287 13209 11299 13243
rect 11241 13203 11299 13209
rect 3016 13144 6500 13172
rect 3016 13132 3022 13144
rect 6546 13132 6552 13184
rect 6604 13132 6610 13184
rect 7009 13175 7067 13181
rect 7009 13141 7021 13175
rect 7055 13172 7067 13175
rect 8018 13172 8024 13184
rect 7055 13144 8024 13172
rect 7055 13141 7067 13144
rect 7009 13135 7067 13141
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 8570 13132 8576 13184
rect 8628 13132 8634 13184
rect 9490 13132 9496 13184
rect 9548 13132 9554 13184
rect 9582 13132 9588 13184
rect 9640 13132 9646 13184
rect 10873 13175 10931 13181
rect 10873 13141 10885 13175
rect 10919 13172 10931 13175
rect 11256 13172 11284 13203
rect 12250 13200 12256 13252
rect 12308 13200 12314 13252
rect 10919 13144 11284 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 12710 13132 12716 13184
rect 12768 13132 12774 13184
rect 13556 13181 13584 13280
rect 13817 13277 13829 13280
rect 13863 13277 13875 13311
rect 13817 13271 13875 13277
rect 13722 13200 13728 13252
rect 13780 13240 13786 13252
rect 14642 13240 14648 13252
rect 13780 13212 14648 13240
rect 13780 13200 13786 13212
rect 14642 13200 14648 13212
rect 14700 13240 14706 13252
rect 15013 13243 15071 13249
rect 15013 13240 15025 13243
rect 14700 13212 15025 13240
rect 14700 13200 14706 13212
rect 15013 13209 15025 13212
rect 15059 13209 15071 13243
rect 15013 13203 15071 13209
rect 15194 13200 15200 13252
rect 15252 13200 15258 13252
rect 16666 13200 16672 13252
rect 16724 13200 16730 13252
rect 13541 13175 13599 13181
rect 13541 13141 13553 13175
rect 13587 13141 13599 13175
rect 13541 13135 13599 13141
rect 13630 13132 13636 13184
rect 13688 13132 13694 13184
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 15286 13172 15292 13184
rect 13872 13144 15292 13172
rect 13872 13132 13878 13144
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 15562 13132 15568 13184
rect 15620 13172 15626 13184
rect 16485 13175 16543 13181
rect 16485 13172 16497 13175
rect 15620 13144 16497 13172
rect 15620 13132 15626 13144
rect 16485 13141 16497 13144
rect 16531 13141 16543 13175
rect 16776 13172 16804 13348
rect 16868 13308 16896 13404
rect 17773 13311 17831 13317
rect 17773 13308 17785 13311
rect 16868 13280 17785 13308
rect 17773 13277 17785 13280
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 16853 13243 16911 13249
rect 16853 13209 16865 13243
rect 16899 13240 16911 13243
rect 17880 13240 17908 13472
rect 16899 13212 17908 13240
rect 18233 13243 18291 13249
rect 16899 13209 16911 13212
rect 16853 13203 16911 13209
rect 18233 13209 18245 13243
rect 18279 13240 18291 13243
rect 18322 13240 18328 13252
rect 18279 13212 18328 13240
rect 18279 13209 18291 13212
rect 18233 13203 18291 13209
rect 18322 13200 18328 13212
rect 18380 13200 18386 13252
rect 18433 13175 18491 13181
rect 18433 13172 18445 13175
rect 16776 13144 18445 13172
rect 16485 13135 16543 13141
rect 18433 13141 18445 13144
rect 18479 13172 18491 13175
rect 18524 13172 18552 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 19702 13472 19708 13524
rect 19760 13472 19766 13524
rect 20622 13512 20628 13524
rect 19996 13484 20628 13512
rect 18601 13447 18659 13453
rect 18601 13413 18613 13447
rect 18647 13444 18659 13447
rect 19334 13444 19340 13456
rect 18647 13416 19340 13444
rect 18647 13413 18659 13416
rect 18601 13407 18659 13413
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 18690 13268 18696 13320
rect 18748 13308 18754 13320
rect 18748 13283 18888 13308
rect 18748 13280 18889 13283
rect 18748 13268 18754 13280
rect 18831 13277 18889 13280
rect 18831 13243 18843 13277
rect 18877 13243 18889 13277
rect 19610 13268 19616 13320
rect 19668 13308 19674 13320
rect 19996 13317 20024 13484
rect 20622 13472 20628 13484
rect 20680 13472 20686 13524
rect 27433 13515 27491 13521
rect 24412 13484 27108 13512
rect 20438 13444 20444 13456
rect 20088 13416 20444 13444
rect 20088 13320 20116 13416
rect 20438 13404 20444 13416
rect 20496 13404 20502 13456
rect 20809 13447 20867 13453
rect 20809 13413 20821 13447
rect 20855 13444 20867 13447
rect 21818 13444 21824 13456
rect 20855 13416 21824 13444
rect 20855 13413 20867 13416
rect 20809 13407 20867 13413
rect 21818 13404 21824 13416
rect 21876 13404 21882 13456
rect 22649 13447 22707 13453
rect 22649 13413 22661 13447
rect 22695 13444 22707 13447
rect 22738 13444 22744 13456
rect 22695 13416 22744 13444
rect 22695 13413 22707 13416
rect 22649 13407 22707 13413
rect 22738 13404 22744 13416
rect 22796 13404 22802 13456
rect 22922 13404 22928 13456
rect 22980 13444 22986 13456
rect 23842 13444 23848 13456
rect 22980 13416 23848 13444
rect 22980 13404 22986 13416
rect 23842 13404 23848 13416
rect 23900 13404 23906 13456
rect 24412 13376 24440 13484
rect 26970 13444 26976 13456
rect 20180 13348 20576 13376
rect 19981 13311 20039 13317
rect 19981 13308 19993 13311
rect 19668 13280 19993 13308
rect 19668 13268 19674 13280
rect 19981 13277 19993 13280
rect 20027 13277 20039 13311
rect 19981 13271 20039 13277
rect 20070 13268 20076 13320
rect 20128 13268 20134 13320
rect 20180 13317 20208 13348
rect 20548 13320 20576 13348
rect 21008 13348 24440 13376
rect 24504 13416 26976 13444
rect 20165 13311 20223 13317
rect 20165 13277 20177 13311
rect 20211 13277 20223 13311
rect 20165 13271 20223 13277
rect 20349 13311 20407 13317
rect 20349 13277 20361 13311
rect 20395 13277 20407 13311
rect 20349 13271 20407 13277
rect 18831 13237 18889 13243
rect 19061 13243 19119 13249
rect 19061 13209 19073 13243
rect 19107 13240 19119 13243
rect 19150 13240 19156 13252
rect 19107 13212 19156 13240
rect 19107 13209 19119 13212
rect 19061 13203 19119 13209
rect 19150 13200 19156 13212
rect 19208 13200 19214 13252
rect 20364 13240 20392 13271
rect 20530 13268 20536 13320
rect 20588 13268 20594 13320
rect 20441 13243 20499 13249
rect 20441 13240 20453 13243
rect 20180 13212 20453 13240
rect 20180 13184 20208 13212
rect 20441 13209 20453 13212
rect 20487 13209 20499 13243
rect 20548 13240 20576 13268
rect 21008 13249 21036 13348
rect 21082 13268 21088 13320
rect 21140 13268 21146 13320
rect 21358 13268 21364 13320
rect 21416 13268 21422 13320
rect 21726 13268 21732 13320
rect 21784 13268 21790 13320
rect 22370 13268 22376 13320
rect 22428 13268 22434 13320
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13308 22615 13311
rect 22925 13311 22983 13317
rect 22925 13308 22937 13311
rect 22603 13280 22937 13308
rect 22603 13277 22615 13280
rect 22557 13271 22615 13277
rect 22925 13277 22937 13280
rect 22971 13277 22983 13311
rect 22925 13271 22983 13277
rect 20641 13243 20699 13249
rect 20641 13240 20653 13243
rect 20548 13212 20653 13240
rect 20441 13203 20499 13209
rect 20641 13209 20653 13212
rect 20687 13209 20699 13243
rect 20641 13203 20699 13209
rect 20993 13243 21051 13249
rect 20993 13209 21005 13243
rect 21039 13209 21051 13243
rect 22572 13240 22600 13271
rect 20993 13203 21051 13209
rect 21192 13212 22600 13240
rect 22940 13240 22968 13271
rect 23198 13268 23204 13320
rect 23256 13308 23262 13320
rect 23477 13311 23535 13317
rect 23477 13308 23489 13311
rect 23256 13280 23489 13308
rect 23256 13268 23262 13280
rect 23477 13277 23489 13280
rect 23523 13277 23535 13311
rect 23477 13271 23535 13277
rect 24118 13268 24124 13320
rect 24176 13308 24182 13320
rect 24397 13311 24455 13317
rect 24397 13308 24409 13311
rect 24176 13280 24409 13308
rect 24176 13268 24182 13280
rect 24397 13277 24409 13280
rect 24443 13277 24455 13311
rect 24397 13271 24455 13277
rect 24504 13252 24532 13416
rect 25774 13336 25780 13388
rect 25832 13376 25838 13388
rect 26234 13376 26240 13388
rect 25832 13348 26004 13376
rect 25832 13336 25838 13348
rect 24673 13311 24731 13317
rect 24673 13277 24685 13311
rect 24719 13308 24731 13311
rect 24854 13308 24860 13320
rect 24719 13280 24860 13308
rect 24719 13277 24731 13280
rect 24673 13271 24731 13277
rect 24854 13268 24860 13280
rect 24912 13268 24918 13320
rect 25590 13268 25596 13320
rect 25648 13308 25654 13320
rect 25685 13311 25743 13317
rect 25685 13308 25697 13311
rect 25648 13280 25697 13308
rect 25648 13268 25654 13280
rect 25685 13277 25697 13280
rect 25731 13277 25743 13311
rect 25685 13271 25743 13277
rect 25866 13268 25872 13320
rect 25924 13268 25930 13320
rect 25976 13317 26004 13348
rect 26068 13348 26240 13376
rect 25961 13311 26019 13317
rect 25961 13277 25973 13311
rect 26007 13277 26019 13311
rect 25961 13271 26019 13277
rect 23293 13243 23351 13249
rect 23293 13240 23305 13243
rect 22940 13212 23305 13240
rect 18479 13144 18552 13172
rect 18479 13141 18491 13144
rect 18433 13135 18491 13141
rect 18690 13132 18696 13184
rect 18748 13132 18754 13184
rect 20162 13132 20168 13184
rect 20220 13132 20226 13184
rect 20530 13132 20536 13184
rect 20588 13172 20594 13184
rect 21008 13172 21036 13203
rect 21192 13184 21220 13212
rect 23293 13209 23305 13212
rect 23339 13209 23351 13243
rect 23293 13203 23351 13209
rect 23661 13243 23719 13249
rect 23661 13209 23673 13243
rect 23707 13240 23719 13243
rect 24486 13240 24492 13252
rect 23707 13212 24492 13240
rect 23707 13209 23719 13212
rect 23661 13203 23719 13209
rect 24486 13200 24492 13212
rect 24544 13200 24550 13252
rect 24765 13243 24823 13249
rect 24765 13209 24777 13243
rect 24811 13240 24823 13243
rect 25498 13240 25504 13252
rect 24811 13212 25504 13240
rect 24811 13209 24823 13212
rect 24765 13203 24823 13209
rect 25498 13200 25504 13212
rect 25556 13200 25562 13252
rect 26068 13240 26096 13348
rect 26234 13336 26240 13348
rect 26292 13336 26298 13388
rect 26344 13385 26372 13416
rect 26970 13404 26976 13416
rect 27028 13404 27034 13456
rect 27080 13444 27108 13484
rect 27433 13481 27445 13515
rect 27479 13512 27491 13515
rect 27798 13512 27804 13524
rect 27479 13484 27804 13512
rect 27479 13481 27491 13484
rect 27433 13475 27491 13481
rect 27798 13472 27804 13484
rect 27856 13472 27862 13524
rect 28077 13515 28135 13521
rect 28077 13481 28089 13515
rect 28123 13512 28135 13515
rect 28166 13512 28172 13524
rect 28123 13484 28172 13512
rect 28123 13481 28135 13484
rect 28077 13475 28135 13481
rect 28166 13472 28172 13484
rect 28224 13472 28230 13524
rect 28994 13472 29000 13524
rect 29052 13512 29058 13524
rect 29089 13515 29147 13521
rect 29089 13512 29101 13515
rect 29052 13484 29101 13512
rect 29052 13472 29058 13484
rect 29089 13481 29101 13484
rect 29135 13481 29147 13515
rect 29089 13475 29147 13481
rect 29178 13472 29184 13524
rect 29236 13512 29242 13524
rect 29236 13484 30328 13512
rect 29236 13472 29242 13484
rect 30300 13456 30328 13484
rect 32398 13472 32404 13524
rect 32456 13512 32462 13524
rect 33137 13515 33195 13521
rect 33137 13512 33149 13515
rect 32456 13484 33149 13512
rect 32456 13472 32462 13484
rect 33137 13481 33149 13484
rect 33183 13481 33195 13515
rect 33137 13475 33195 13481
rect 33226 13472 33232 13524
rect 33284 13472 33290 13524
rect 33410 13472 33416 13524
rect 33468 13512 33474 13524
rect 33689 13515 33747 13521
rect 33689 13512 33701 13515
rect 33468 13484 33701 13512
rect 33468 13472 33474 13484
rect 33689 13481 33701 13484
rect 33735 13481 33747 13515
rect 33689 13475 33747 13481
rect 28261 13447 28319 13453
rect 28261 13444 28273 13447
rect 27080 13416 28273 13444
rect 28261 13413 28273 13416
rect 28307 13444 28319 13447
rect 28350 13444 28356 13456
rect 28307 13416 28356 13444
rect 28307 13413 28319 13416
rect 28261 13407 28319 13413
rect 28350 13404 28356 13416
rect 28408 13404 28414 13456
rect 30282 13404 30288 13456
rect 30340 13404 30346 13456
rect 31202 13404 31208 13456
rect 31260 13444 31266 13456
rect 32122 13444 32128 13456
rect 31260 13416 32128 13444
rect 31260 13404 31266 13416
rect 32122 13404 32128 13416
rect 32180 13404 32186 13456
rect 33428 13444 33456 13472
rect 32968 13416 33456 13444
rect 32968 13385 32996 13416
rect 26329 13379 26387 13385
rect 26329 13345 26341 13379
rect 26375 13345 26387 13379
rect 26329 13339 26387 13345
rect 26697 13379 26755 13385
rect 26697 13345 26709 13379
rect 26743 13376 26755 13379
rect 28997 13379 29055 13385
rect 28997 13376 29009 13379
rect 26743 13348 27016 13376
rect 26743 13345 26755 13348
rect 26697 13339 26755 13345
rect 26145 13311 26203 13317
rect 26145 13277 26157 13311
rect 26191 13277 26203 13311
rect 26145 13271 26203 13277
rect 25700 13212 26096 13240
rect 26160 13240 26188 13271
rect 26510 13268 26516 13320
rect 26568 13268 26574 13320
rect 26786 13268 26792 13320
rect 26844 13268 26850 13320
rect 26988 13317 27016 13348
rect 27448 13348 29009 13376
rect 26973 13311 27031 13317
rect 26973 13277 26985 13311
rect 27019 13277 27031 13311
rect 26973 13271 27031 13277
rect 27062 13268 27068 13320
rect 27120 13268 27126 13320
rect 27154 13268 27160 13320
rect 27212 13308 27218 13320
rect 27448 13308 27476 13348
rect 28997 13345 29009 13348
rect 29043 13345 29055 13379
rect 32953 13379 33011 13385
rect 28997 13339 29055 13345
rect 29196 13348 29776 13376
rect 27212 13280 27476 13308
rect 28353 13311 28411 13317
rect 27212 13268 27218 13280
rect 28353 13277 28365 13311
rect 28399 13277 28411 13311
rect 28353 13271 28411 13277
rect 28445 13311 28503 13317
rect 28445 13277 28457 13311
rect 28491 13277 28503 13311
rect 28445 13271 28503 13277
rect 26694 13240 26700 13252
rect 26160 13212 26700 13240
rect 20588 13144 21036 13172
rect 20588 13132 20594 13144
rect 21174 13132 21180 13184
rect 21232 13132 21238 13184
rect 21542 13132 21548 13184
rect 21600 13132 21606 13184
rect 22186 13132 22192 13184
rect 22244 13172 22250 13184
rect 25700 13172 25728 13212
rect 26694 13200 26700 13212
rect 26752 13200 26758 13252
rect 22244 13144 25728 13172
rect 22244 13132 22250 13144
rect 25774 13132 25780 13184
rect 25832 13132 25838 13184
rect 26510 13132 26516 13184
rect 26568 13172 26574 13184
rect 27172 13172 27200 13268
rect 26568 13144 27200 13172
rect 28368 13172 28396 13271
rect 28460 13240 28488 13271
rect 28534 13268 28540 13320
rect 28592 13268 28598 13320
rect 28721 13311 28779 13317
rect 28721 13277 28733 13311
rect 28767 13308 28779 13311
rect 29196 13308 29224 13348
rect 28767 13280 29224 13308
rect 28767 13277 28779 13280
rect 28721 13271 28779 13277
rect 29270 13268 29276 13320
rect 29328 13268 29334 13320
rect 29454 13268 29460 13320
rect 29512 13308 29518 13320
rect 29748 13317 29776 13348
rect 32953 13345 32965 13379
rect 32999 13345 33011 13379
rect 34057 13379 34115 13385
rect 34057 13376 34069 13379
rect 32953 13339 33011 13345
rect 33152 13348 34069 13376
rect 33152 13320 33180 13348
rect 34057 13345 34069 13348
rect 34103 13345 34115 13379
rect 34057 13339 34115 13345
rect 29549 13311 29607 13317
rect 29549 13308 29561 13311
rect 29512 13280 29561 13308
rect 29512 13268 29518 13280
rect 29549 13277 29561 13280
rect 29595 13277 29607 13311
rect 29549 13271 29607 13277
rect 29733 13311 29791 13317
rect 29733 13277 29745 13311
rect 29779 13308 29791 13311
rect 31202 13308 31208 13320
rect 29779 13280 31208 13308
rect 29779 13277 29791 13280
rect 29733 13271 29791 13277
rect 31202 13268 31208 13280
rect 31260 13268 31266 13320
rect 32858 13268 32864 13320
rect 32916 13268 32922 13320
rect 33134 13268 33140 13320
rect 33192 13268 33198 13320
rect 33413 13311 33471 13317
rect 33413 13277 33425 13311
rect 33459 13277 33471 13311
rect 33413 13271 33471 13277
rect 28460 13212 29684 13240
rect 29656 13184 29684 13212
rect 31294 13200 31300 13252
rect 31352 13240 31358 13252
rect 31662 13240 31668 13252
rect 31352 13212 31668 13240
rect 31352 13200 31358 13212
rect 31662 13200 31668 13212
rect 31720 13240 31726 13252
rect 32493 13243 32551 13249
rect 32493 13240 32505 13243
rect 31720 13212 32505 13240
rect 31720 13200 31726 13212
rect 32493 13209 32505 13212
rect 32539 13209 32551 13243
rect 32493 13203 32551 13209
rect 32582 13200 32588 13252
rect 32640 13200 32646 13252
rect 33428 13240 33456 13271
rect 33502 13268 33508 13320
rect 33560 13268 33566 13320
rect 33870 13268 33876 13320
rect 33928 13268 33934 13320
rect 32968 13212 33456 13240
rect 32968 13184 32996 13212
rect 28442 13172 28448 13184
rect 28368 13144 28448 13172
rect 26568 13132 26574 13144
rect 28442 13132 28448 13144
rect 28500 13172 28506 13184
rect 28902 13172 28908 13184
rect 28500 13144 28908 13172
rect 28500 13132 28506 13144
rect 28902 13132 28908 13144
rect 28960 13132 28966 13184
rect 29638 13132 29644 13184
rect 29696 13132 29702 13184
rect 32950 13132 32956 13184
rect 33008 13132 33014 13184
rect 1104 13082 38272 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38272 13082
rect 1104 13008 38272 13030
rect 3145 12971 3203 12977
rect 3145 12937 3157 12971
rect 3191 12968 3203 12971
rect 3970 12968 3976 12980
rect 3191 12940 3976 12968
rect 3191 12937 3203 12940
rect 3145 12931 3203 12937
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 4614 12928 4620 12980
rect 4672 12968 4678 12980
rect 4985 12971 5043 12977
rect 4985 12968 4997 12971
rect 4672 12940 4997 12968
rect 4672 12928 4678 12940
rect 4985 12937 4997 12940
rect 5031 12937 5043 12971
rect 4985 12931 5043 12937
rect 6546 12928 6552 12980
rect 6604 12928 6610 12980
rect 7024 12940 7788 12968
rect 4065 12903 4123 12909
rect 4065 12869 4077 12903
rect 4111 12900 4123 12903
rect 4525 12903 4583 12909
rect 4525 12900 4537 12903
rect 4111 12872 4537 12900
rect 4111 12869 4123 12872
rect 4065 12863 4123 12869
rect 4525 12869 4537 12872
rect 4571 12869 4583 12903
rect 6564 12900 6592 12928
rect 4525 12863 4583 12869
rect 6012 12872 6592 12900
rect 1394 12792 1400 12844
rect 1452 12792 1458 12844
rect 2958 12832 2964 12844
rect 2806 12804 2964 12832
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3970 12792 3976 12844
rect 4028 12792 4034 12844
rect 4430 12792 4436 12844
rect 4488 12792 4494 12844
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4706 12832 4712 12844
rect 4663 12804 4712 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 1670 12724 1676 12776
rect 1728 12724 1734 12776
rect 3878 12724 3884 12776
rect 3936 12764 3942 12776
rect 4157 12767 4215 12773
rect 4157 12764 4169 12767
rect 3936 12736 4169 12764
rect 3936 12724 3942 12736
rect 4157 12733 4169 12736
rect 4203 12733 4215 12767
rect 4157 12727 4215 12733
rect 3786 12656 3792 12708
rect 3844 12696 3850 12708
rect 4632 12696 4660 12795
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12832 5227 12835
rect 5810 12832 5816 12844
rect 5215 12804 5816 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 6012 12841 6040 12872
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 7024 12900 7052 12940
rect 6972 12872 7130 12900
rect 6972 12860 6978 12872
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6362 12792 6368 12844
rect 6420 12792 6426 12844
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6196 12736 6653 12764
rect 6196 12705 6224 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 7760 12764 7788 12940
rect 8018 12928 8024 12980
rect 8076 12968 8082 12980
rect 8113 12971 8171 12977
rect 8113 12968 8125 12971
rect 8076 12940 8125 12968
rect 8076 12928 8082 12940
rect 8113 12937 8125 12940
rect 8159 12937 8171 12971
rect 9858 12968 9864 12980
rect 8113 12931 8171 12937
rect 8312 12940 9864 12968
rect 8312 12841 8340 12940
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 10410 12928 10416 12980
rect 10468 12928 10474 12980
rect 13630 12928 13636 12980
rect 13688 12928 13694 12980
rect 13814 12928 13820 12980
rect 13872 12928 13878 12980
rect 14921 12971 14979 12977
rect 14921 12937 14933 12971
rect 14967 12968 14979 12971
rect 15194 12968 15200 12980
rect 14967 12940 15200 12968
rect 14967 12937 14979 12940
rect 14921 12931 14979 12937
rect 15194 12928 15200 12940
rect 15252 12928 15258 12980
rect 19731 12971 19789 12977
rect 19731 12937 19743 12971
rect 19777 12968 19789 12971
rect 20070 12968 20076 12980
rect 19777 12940 20076 12968
rect 19777 12937 19789 12940
rect 19731 12931 19789 12937
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 20349 12971 20407 12977
rect 20349 12937 20361 12971
rect 20395 12968 20407 12971
rect 21174 12968 21180 12980
rect 20395 12940 21180 12968
rect 20395 12937 20407 12940
rect 20349 12931 20407 12937
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 21637 12971 21695 12977
rect 21637 12937 21649 12971
rect 21683 12968 21695 12971
rect 21726 12968 21732 12980
rect 21683 12940 21732 12968
rect 21683 12937 21695 12940
rect 21637 12931 21695 12937
rect 21726 12928 21732 12940
rect 21784 12928 21790 12980
rect 22066 12940 23243 12968
rect 8570 12860 8576 12912
rect 8628 12860 8634 12912
rect 10428 12900 10456 12928
rect 13449 12903 13507 12909
rect 10428 12872 10640 12900
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 9674 12792 9680 12844
rect 9732 12792 9738 12844
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10612 12841 10640 12872
rect 13449 12869 13461 12903
rect 13495 12900 13507 12903
rect 13648 12900 13676 12928
rect 13495 12872 13676 12900
rect 13832 12900 13860 12928
rect 13832 12872 13938 12900
rect 13495 12869 13507 12872
rect 13449 12863 13507 12869
rect 19242 12860 19248 12912
rect 19300 12900 19306 12912
rect 19521 12903 19579 12909
rect 19521 12900 19533 12903
rect 19300 12872 19533 12900
rect 19300 12860 19306 12872
rect 19521 12869 19533 12872
rect 19567 12869 19579 12903
rect 20088 12900 20116 12928
rect 20088 12872 20576 12900
rect 19521 12863 19579 12869
rect 10321 12835 10379 12841
rect 10321 12832 10333 12835
rect 10284 12804 10333 12832
rect 10284 12792 10290 12804
rect 10321 12801 10333 12804
rect 10367 12801 10379 12835
rect 10505 12835 10563 12841
rect 10505 12832 10517 12835
rect 10321 12795 10379 12801
rect 10428 12804 10517 12832
rect 9692 12764 9720 12792
rect 7760 12736 9720 12764
rect 6641 12727 6699 12733
rect 3844 12668 4660 12696
rect 6181 12699 6239 12705
rect 3844 12656 3850 12668
rect 6181 12665 6193 12699
rect 6227 12665 6239 12699
rect 6181 12659 6239 12665
rect 9582 12656 9588 12708
rect 9640 12696 9646 12708
rect 10045 12699 10103 12705
rect 10045 12696 10057 12699
rect 9640 12668 10057 12696
rect 9640 12656 9646 12668
rect 10045 12665 10057 12668
rect 10091 12696 10103 12699
rect 10428 12696 10456 12804
rect 10505 12801 10517 12804
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 10597 12835 10655 12841
rect 10597 12801 10609 12835
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 11940 12804 12664 12832
rect 11940 12792 11946 12804
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 12032 12736 12265 12764
rect 12032 12724 12038 12736
rect 12253 12733 12265 12736
rect 12299 12733 12311 12767
rect 12636 12764 12664 12804
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 13081 12835 13139 12841
rect 13081 12832 13093 12835
rect 12768 12804 13093 12832
rect 12768 12792 12774 12804
rect 13081 12801 13093 12804
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 14918 12792 14924 12844
rect 14976 12792 14982 12844
rect 15470 12792 15476 12844
rect 15528 12792 15534 12844
rect 15580 12804 16804 12832
rect 13170 12764 13176 12776
rect 12636 12736 13176 12764
rect 12253 12727 12311 12733
rect 13170 12724 13176 12736
rect 13228 12724 13234 12776
rect 14936 12764 14964 12792
rect 15580 12773 15608 12804
rect 15565 12767 15623 12773
rect 15565 12764 15577 12767
rect 14936 12736 15577 12764
rect 15565 12733 15577 12736
rect 15611 12733 15623 12767
rect 15565 12727 15623 12733
rect 15654 12724 15660 12776
rect 15712 12724 15718 12776
rect 16776 12764 16804 12804
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 19536 12832 19564 12863
rect 20162 12832 20168 12844
rect 19536 12804 20168 12832
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 20548 12841 20576 12872
rect 20990 12860 20996 12912
rect 21048 12900 21054 12912
rect 21542 12900 21548 12912
rect 21048 12872 21548 12900
rect 21048 12860 21054 12872
rect 21542 12860 21548 12872
rect 21600 12900 21606 12912
rect 22066 12900 22094 12940
rect 21600 12872 22094 12900
rect 23215 12900 23243 12940
rect 24762 12928 24768 12980
rect 24820 12968 24826 12980
rect 24857 12971 24915 12977
rect 24857 12968 24869 12971
rect 24820 12940 24869 12968
rect 24820 12928 24826 12940
rect 24857 12937 24869 12940
rect 24903 12937 24915 12971
rect 24857 12931 24915 12937
rect 25866 12928 25872 12980
rect 25924 12968 25930 12980
rect 26237 12971 26295 12977
rect 26237 12968 26249 12971
rect 25924 12940 26249 12968
rect 25924 12928 25930 12940
rect 26237 12937 26249 12940
rect 26283 12937 26295 12971
rect 26237 12931 26295 12937
rect 26694 12928 26700 12980
rect 26752 12928 26758 12980
rect 29638 12928 29644 12980
rect 29696 12928 29702 12980
rect 31202 12928 31208 12980
rect 31260 12968 31266 12980
rect 31260 12940 31524 12968
rect 31260 12928 31266 12940
rect 26712 12900 26740 12928
rect 23215 12872 24992 12900
rect 21600 12860 21606 12872
rect 20533 12835 20591 12841
rect 20533 12801 20545 12835
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 17589 12767 17647 12773
rect 17589 12764 17601 12767
rect 16776 12736 17601 12764
rect 17589 12733 17601 12736
rect 17635 12764 17647 12767
rect 19978 12764 19984 12776
rect 17635 12736 19984 12764
rect 17635 12733 17647 12736
rect 17589 12727 17647 12733
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 21100 12764 21128 12795
rect 21450 12792 21456 12844
rect 21508 12792 21514 12844
rect 21818 12792 21824 12844
rect 21876 12792 21882 12844
rect 23198 12832 23204 12844
rect 22066 12804 23204 12832
rect 21836 12764 21864 12792
rect 21100 12736 21864 12764
rect 10091 12668 10456 12696
rect 14476 12668 16436 12696
rect 10091 12665 10103 12668
rect 10045 12659 10103 12665
rect 3050 12588 3056 12640
rect 3108 12628 3114 12640
rect 3605 12631 3663 12637
rect 3605 12628 3617 12631
rect 3108 12600 3617 12628
rect 3108 12588 3114 12600
rect 3605 12597 3617 12600
rect 3651 12597 3663 12631
rect 3605 12591 3663 12597
rect 10134 12588 10140 12640
rect 10192 12588 10198 12640
rect 10244 12628 10272 12668
rect 14476 12628 14504 12668
rect 16408 12640 16436 12668
rect 10244 12600 14504 12628
rect 15102 12588 15108 12640
rect 15160 12588 15166 12640
rect 16390 12588 16396 12640
rect 16448 12588 16454 12640
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 19705 12631 19763 12637
rect 19705 12628 19717 12631
rect 19484 12600 19717 12628
rect 19484 12588 19490 12600
rect 19705 12597 19717 12600
rect 19751 12597 19763 12631
rect 19705 12591 19763 12597
rect 19886 12588 19892 12640
rect 19944 12588 19950 12640
rect 20165 12631 20223 12637
rect 20165 12597 20177 12631
rect 20211 12628 20223 12631
rect 20622 12628 20628 12640
rect 20211 12600 20628 12628
rect 20211 12597 20223 12600
rect 20165 12591 20223 12597
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 21358 12588 21364 12640
rect 21416 12628 21422 12640
rect 21453 12631 21511 12637
rect 21453 12628 21465 12631
rect 21416 12600 21465 12628
rect 21416 12588 21422 12600
rect 21453 12597 21465 12600
rect 21499 12628 21511 12631
rect 22066 12628 22094 12804
rect 22186 12724 22192 12776
rect 22244 12724 22250 12776
rect 22278 12724 22284 12776
rect 22336 12724 22342 12776
rect 22388 12773 22416 12804
rect 23198 12792 23204 12804
rect 23256 12792 23262 12844
rect 24210 12792 24216 12844
rect 24268 12832 24274 12844
rect 24964 12841 24992 12872
rect 26344 12872 26648 12900
rect 26712 12872 26832 12900
rect 26344 12844 26372 12872
rect 24949 12835 25007 12841
rect 24268 12804 24716 12832
rect 24268 12792 24274 12804
rect 22373 12767 22431 12773
rect 22373 12733 22385 12767
rect 22419 12733 22431 12767
rect 22373 12727 22431 12733
rect 24118 12724 24124 12776
rect 24176 12724 24182 12776
rect 24302 12724 24308 12776
rect 24360 12764 24366 12776
rect 24397 12767 24455 12773
rect 24397 12764 24409 12767
rect 24360 12736 24409 12764
rect 24360 12724 24366 12736
rect 24397 12733 24409 12736
rect 24443 12733 24455 12767
rect 24397 12727 24455 12733
rect 24486 12724 24492 12776
rect 24544 12724 24550 12776
rect 24688 12773 24716 12804
rect 24949 12801 24961 12835
rect 24995 12801 25007 12835
rect 24949 12795 25007 12801
rect 25041 12835 25099 12841
rect 25041 12801 25053 12835
rect 25087 12832 25099 12835
rect 25590 12832 25596 12844
rect 25087 12804 25596 12832
rect 25087 12801 25099 12804
rect 25041 12795 25099 12801
rect 25590 12792 25596 12804
rect 25648 12792 25654 12844
rect 26326 12792 26332 12844
rect 26384 12792 26390 12844
rect 26421 12835 26479 12841
rect 26421 12801 26433 12835
rect 26467 12801 26479 12835
rect 26421 12795 26479 12801
rect 24581 12767 24639 12773
rect 24581 12733 24593 12767
rect 24627 12733 24639 12767
rect 24581 12727 24639 12733
rect 24673 12767 24731 12773
rect 24673 12733 24685 12767
rect 24719 12733 24731 12767
rect 24673 12727 24731 12733
rect 22302 12696 22330 12724
rect 22554 12696 22560 12708
rect 22302 12668 22560 12696
rect 22554 12656 22560 12668
rect 22612 12696 22618 12708
rect 24136 12696 24164 12724
rect 24596 12696 24624 12727
rect 25222 12724 25228 12776
rect 25280 12724 25286 12776
rect 26436 12764 26464 12795
rect 26510 12792 26516 12844
rect 26568 12792 26574 12844
rect 26620 12832 26648 12872
rect 26804 12841 26832 12872
rect 26697 12835 26755 12841
rect 26697 12832 26709 12835
rect 26620 12804 26709 12832
rect 26697 12801 26709 12804
rect 26743 12801 26755 12835
rect 26697 12795 26755 12801
rect 26789 12835 26847 12841
rect 26789 12801 26801 12835
rect 26835 12801 26847 12835
rect 26789 12795 26847 12801
rect 29089 12835 29147 12841
rect 29089 12801 29101 12835
rect 29135 12832 29147 12835
rect 29656 12832 29684 12928
rect 31496 12909 31524 12940
rect 31846 12928 31852 12980
rect 31904 12928 31910 12980
rect 32858 12928 32864 12980
rect 32916 12928 32922 12980
rect 33134 12928 33140 12980
rect 33192 12928 33198 12980
rect 31481 12903 31539 12909
rect 29135 12804 29684 12832
rect 29748 12872 31340 12900
rect 29135 12801 29147 12804
rect 29089 12795 29147 12801
rect 26878 12764 26884 12776
rect 26436 12736 26884 12764
rect 26878 12724 26884 12736
rect 26936 12724 26942 12776
rect 28166 12724 28172 12776
rect 28224 12764 28230 12776
rect 29365 12767 29423 12773
rect 29365 12764 29377 12767
rect 28224 12736 29377 12764
rect 28224 12724 28230 12736
rect 29365 12733 29377 12736
rect 29411 12764 29423 12767
rect 29748 12764 29776 12872
rect 30006 12792 30012 12844
rect 30064 12792 30070 12844
rect 30374 12792 30380 12844
rect 30432 12832 30438 12844
rect 30650 12832 30656 12844
rect 30432 12804 30656 12832
rect 30432 12792 30438 12804
rect 30650 12792 30656 12804
rect 30708 12792 30714 12844
rect 31202 12792 31208 12844
rect 31260 12792 31266 12844
rect 29411 12736 29776 12764
rect 29411 12733 29423 12736
rect 29365 12727 29423 12733
rect 24854 12696 24860 12708
rect 22612 12668 24860 12696
rect 22612 12656 22618 12668
rect 24854 12656 24860 12668
rect 24912 12656 24918 12708
rect 25774 12656 25780 12708
rect 25832 12696 25838 12708
rect 28994 12696 29000 12708
rect 25832 12668 29000 12696
rect 25832 12656 25838 12668
rect 28994 12656 29000 12668
rect 29052 12656 29058 12708
rect 29086 12656 29092 12708
rect 29144 12696 29150 12708
rect 29181 12699 29239 12705
rect 29181 12696 29193 12699
rect 29144 12668 29193 12696
rect 29144 12656 29150 12668
rect 29181 12665 29193 12668
rect 29227 12696 29239 12699
rect 30024 12696 30052 12792
rect 30282 12724 30288 12776
rect 30340 12764 30346 12776
rect 30561 12767 30619 12773
rect 30561 12764 30573 12767
rect 30340 12736 30573 12764
rect 30340 12724 30346 12736
rect 30561 12733 30573 12736
rect 30607 12733 30619 12767
rect 30561 12727 30619 12733
rect 29227 12668 30052 12696
rect 31021 12699 31079 12705
rect 29227 12665 29239 12668
rect 29181 12659 29239 12665
rect 31021 12665 31033 12699
rect 31067 12696 31079 12699
rect 31220 12696 31248 12792
rect 31312 12764 31340 12872
rect 31481 12869 31493 12903
rect 31527 12869 31539 12903
rect 31481 12863 31539 12869
rect 31697 12903 31755 12909
rect 31697 12869 31709 12903
rect 31743 12900 31755 12903
rect 32493 12903 32551 12909
rect 32493 12900 32505 12903
rect 31743 12872 32505 12900
rect 31743 12869 31755 12872
rect 31697 12863 31755 12869
rect 32493 12869 32505 12872
rect 32539 12869 32551 12903
rect 32493 12863 32551 12869
rect 31386 12792 31392 12844
rect 31444 12832 31450 12844
rect 33152 12841 33180 12928
rect 32125 12835 32183 12841
rect 32125 12832 32137 12835
rect 31444 12804 32137 12832
rect 31444 12792 31450 12804
rect 32125 12801 32137 12804
rect 32171 12801 32183 12835
rect 32125 12795 32183 12801
rect 32309 12835 32367 12841
rect 32309 12801 32321 12835
rect 32355 12801 32367 12835
rect 32309 12795 32367 12801
rect 33137 12835 33195 12841
rect 33137 12801 33149 12835
rect 33183 12801 33195 12835
rect 33137 12795 33195 12801
rect 31312 12736 31616 12764
rect 31067 12668 31248 12696
rect 31067 12665 31079 12668
rect 31021 12659 31079 12665
rect 21499 12600 22094 12628
rect 21499 12597 21511 12600
rect 21453 12591 21511 12597
rect 25130 12588 25136 12640
rect 25188 12588 25194 12640
rect 29273 12631 29331 12637
rect 29273 12597 29285 12631
rect 29319 12628 29331 12631
rect 30006 12628 30012 12640
rect 29319 12600 30012 12628
rect 29319 12597 29331 12600
rect 29273 12591 29331 12597
rect 30006 12588 30012 12600
rect 30064 12588 30070 12640
rect 31588 12628 31616 12736
rect 31662 12724 31668 12776
rect 31720 12764 31726 12776
rect 32324 12764 32352 12795
rect 33870 12792 33876 12844
rect 33928 12792 33934 12844
rect 31720 12736 32352 12764
rect 31720 12724 31726 12736
rect 32674 12724 32680 12776
rect 32732 12764 32738 12776
rect 32861 12767 32919 12773
rect 32861 12764 32873 12767
rect 32732 12736 32873 12764
rect 32732 12724 32738 12736
rect 32861 12733 32873 12736
rect 32907 12733 32919 12767
rect 32861 12727 32919 12733
rect 33045 12767 33103 12773
rect 33045 12733 33057 12767
rect 33091 12764 33103 12767
rect 33318 12764 33324 12776
rect 33091 12736 33324 12764
rect 33091 12733 33103 12736
rect 33045 12727 33103 12733
rect 33318 12724 33324 12736
rect 33376 12764 33382 12776
rect 33888 12764 33916 12792
rect 33376 12736 33916 12764
rect 33376 12724 33382 12736
rect 32030 12656 32036 12708
rect 32088 12696 32094 12708
rect 32692 12696 32720 12724
rect 32088 12668 32720 12696
rect 32088 12656 32094 12668
rect 31665 12631 31723 12637
rect 31665 12628 31677 12631
rect 31588 12600 31677 12628
rect 31665 12597 31677 12600
rect 31711 12597 31723 12631
rect 31665 12591 31723 12597
rect 1104 12538 38272 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38272 12538
rect 1104 12464 38272 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 1949 12427 2007 12433
rect 1949 12424 1961 12427
rect 1728 12396 1961 12424
rect 1728 12384 1734 12396
rect 1949 12393 1961 12396
rect 1995 12393 2007 12427
rect 1949 12387 2007 12393
rect 3786 12384 3792 12436
rect 3844 12384 3850 12436
rect 3973 12427 4031 12433
rect 3973 12393 3985 12427
rect 4019 12424 4031 12427
rect 4062 12424 4068 12436
rect 4019 12396 4068 12424
rect 4019 12393 4031 12396
rect 3973 12387 4031 12393
rect 3988 12356 4016 12387
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4614 12424 4620 12436
rect 4295 12396 4620 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 5810 12384 5816 12436
rect 5868 12424 5874 12436
rect 6457 12427 6515 12433
rect 6457 12424 6469 12427
rect 5868 12396 6469 12424
rect 5868 12384 5874 12396
rect 6457 12393 6469 12396
rect 6503 12393 6515 12427
rect 6457 12387 6515 12393
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 8846 12424 8852 12436
rect 8619 12396 8852 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 11517 12427 11575 12433
rect 11517 12424 11529 12427
rect 11204 12396 11529 12424
rect 11204 12384 11210 12396
rect 11517 12393 11529 12396
rect 11563 12393 11575 12427
rect 11517 12387 11575 12393
rect 14921 12427 14979 12433
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 15362 12427 15420 12433
rect 15362 12424 15374 12427
rect 14967 12396 15374 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15362 12393 15374 12396
rect 15408 12393 15420 12427
rect 15362 12387 15420 12393
rect 16850 12384 16856 12436
rect 16908 12384 16914 12436
rect 18322 12384 18328 12436
rect 18380 12424 18386 12436
rect 19242 12424 19248 12436
rect 18380 12396 19248 12424
rect 18380 12384 18386 12396
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 21729 12427 21787 12433
rect 21729 12393 21741 12427
rect 21775 12424 21787 12427
rect 22370 12424 22376 12436
rect 21775 12396 22376 12424
rect 21775 12393 21787 12396
rect 21729 12387 21787 12393
rect 22370 12384 22376 12396
rect 22428 12384 22434 12436
rect 23566 12424 23572 12436
rect 22848 12396 23572 12424
rect 2976 12328 4016 12356
rect 2976 12229 3004 12328
rect 3050 12248 3056 12300
rect 3108 12248 3114 12300
rect 3234 12248 3240 12300
rect 3292 12248 3298 12300
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 2961 12223 3019 12229
rect 2179 12192 2636 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2608 12093 2636 12192
rect 2961 12189 2973 12223
rect 3007 12189 3019 12223
rect 3988 12220 4016 12328
rect 4080 12328 15056 12356
rect 4080 12300 4108 12328
rect 4062 12248 4068 12300
rect 4120 12248 4126 12300
rect 6270 12248 6276 12300
rect 6328 12288 6334 12300
rect 6917 12291 6975 12297
rect 6917 12288 6929 12291
rect 6328 12260 6929 12288
rect 6328 12248 6334 12260
rect 6917 12257 6929 12260
rect 6963 12257 6975 12291
rect 6917 12251 6975 12257
rect 7101 12291 7159 12297
rect 7101 12257 7113 12291
rect 7147 12288 7159 12291
rect 7282 12288 7288 12300
rect 7147 12260 7288 12288
rect 7147 12257 7159 12260
rect 7101 12251 7159 12257
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 8846 12248 8852 12300
rect 8904 12288 8910 12300
rect 8904 12260 10180 12288
rect 8904 12248 8910 12260
rect 4249 12223 4307 12229
rect 4249 12220 4261 12223
rect 3988 12192 4261 12220
rect 2961 12183 3019 12189
rect 4249 12189 4261 12192
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12220 8263 12223
rect 8294 12220 8300 12232
rect 8251 12192 8300 12220
rect 8251 12189 8263 12192
rect 8205 12183 8263 12189
rect 3142 12112 3148 12164
rect 3200 12152 3206 12164
rect 4157 12155 4215 12161
rect 4157 12152 4169 12155
rect 3200 12124 4169 12152
rect 3200 12112 3206 12124
rect 4157 12121 4169 12124
rect 4203 12152 4215 12155
rect 4433 12155 4491 12161
rect 4433 12152 4445 12155
rect 4203 12124 4445 12152
rect 4203 12121 4215 12124
rect 4157 12115 4215 12121
rect 4433 12121 4445 12124
rect 4479 12121 4491 12155
rect 4433 12115 4491 12121
rect 2593 12087 2651 12093
rect 2593 12053 2605 12087
rect 2639 12053 2651 12087
rect 2593 12047 2651 12053
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 3947 12087 4005 12093
rect 3947 12084 3959 12087
rect 3476 12056 3959 12084
rect 3476 12044 3482 12056
rect 3947 12053 3959 12056
rect 3993 12084 4005 12087
rect 4540 12084 4568 12183
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12220 8447 12223
rect 8754 12220 8760 12232
rect 8435 12192 8760 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8754 12180 8760 12192
rect 8812 12180 8818 12232
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12220 10011 12223
rect 10042 12220 10048 12232
rect 9999 12192 10048 12220
rect 9999 12189 10011 12192
rect 9953 12183 10011 12189
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10152 12229 10180 12260
rect 11974 12248 11980 12300
rect 12032 12248 12038 12300
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12288 12219 12291
rect 12618 12288 12624 12300
rect 12207 12260 12624 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 12618 12248 12624 12260
rect 12676 12248 12682 12300
rect 13170 12248 13176 12300
rect 13228 12288 13234 12300
rect 15028 12288 15056 12328
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 16448 12328 18460 12356
rect 16448 12316 16454 12328
rect 13228 12260 14872 12288
rect 15028 12260 17632 12288
rect 13228 12248 13234 12260
rect 10137 12223 10195 12229
rect 10137 12189 10149 12223
rect 10183 12220 10195 12223
rect 10226 12220 10232 12232
rect 10183 12192 10232 12220
rect 10183 12189 10195 12192
rect 10137 12183 10195 12189
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 14734 12180 14740 12232
rect 14792 12180 14798 12232
rect 14844 12220 14872 12260
rect 15105 12223 15163 12229
rect 15105 12220 15117 12223
rect 14844 12192 15117 12220
rect 15105 12189 15117 12192
rect 15151 12189 15163 12223
rect 15105 12183 15163 12189
rect 16482 12180 16488 12232
rect 16540 12180 16546 12232
rect 6825 12155 6883 12161
rect 6825 12121 6837 12155
rect 6871 12152 6883 12155
rect 7926 12152 7932 12164
rect 6871 12124 7932 12152
rect 6871 12121 6883 12124
rect 6825 12115 6883 12121
rect 7926 12112 7932 12124
rect 7984 12152 7990 12164
rect 8665 12155 8723 12161
rect 7984 12124 8616 12152
rect 7984 12112 7990 12124
rect 3993 12056 4568 12084
rect 3993 12053 4005 12056
rect 3947 12047 4005 12053
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 8021 12087 8079 12093
rect 8021 12084 8033 12087
rect 7892 12056 8033 12084
rect 7892 12044 7898 12056
rect 8021 12053 8033 12056
rect 8067 12053 8079 12087
rect 8588 12084 8616 12124
rect 8665 12121 8677 12155
rect 8711 12152 8723 12155
rect 9490 12152 9496 12164
rect 8711 12124 9496 12152
rect 8711 12121 8723 12124
rect 8665 12115 8723 12121
rect 9490 12112 9496 12124
rect 9548 12152 9554 12164
rect 11885 12155 11943 12161
rect 11885 12152 11897 12155
rect 9548 12124 11897 12152
rect 9548 12112 9554 12124
rect 11885 12121 11897 12124
rect 11931 12121 11943 12155
rect 11885 12115 11943 12121
rect 9769 12087 9827 12093
rect 9769 12084 9781 12087
rect 8588 12056 9781 12084
rect 8021 12047 8079 12053
rect 9769 12053 9781 12056
rect 9815 12084 9827 12087
rect 15286 12084 15292 12096
rect 9815 12056 15292 12084
rect 9815 12053 9827 12056
rect 9769 12047 9827 12053
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 17604 12093 17632 12260
rect 17770 12248 17776 12300
rect 17828 12288 17834 12300
rect 18141 12291 18199 12297
rect 18141 12288 18153 12291
rect 17828 12260 18153 12288
rect 17828 12248 17834 12260
rect 18141 12257 18153 12260
rect 18187 12288 18199 12291
rect 18322 12288 18328 12300
rect 18187 12260 18328 12288
rect 18187 12257 18199 12260
rect 18141 12251 18199 12257
rect 18322 12248 18328 12260
rect 18380 12248 18386 12300
rect 18432 12297 18460 12328
rect 19886 12316 19892 12368
rect 19944 12356 19950 12368
rect 22848 12356 22876 12396
rect 23566 12384 23572 12396
rect 23624 12424 23630 12436
rect 23624 12396 23796 12424
rect 23624 12384 23630 12396
rect 23661 12359 23719 12365
rect 23661 12356 23673 12359
rect 19944 12328 22876 12356
rect 22940 12328 23673 12356
rect 19944 12316 19950 12328
rect 18417 12291 18475 12297
rect 18417 12257 18429 12291
rect 18463 12257 18475 12291
rect 20806 12288 20812 12300
rect 18417 12251 18475 12257
rect 18708 12260 20812 12288
rect 18230 12180 18236 12232
rect 18288 12220 18294 12232
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 18288 12192 18613 12220
rect 18288 12180 18294 12192
rect 18601 12189 18613 12192
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 18049 12155 18107 12161
rect 18049 12121 18061 12155
rect 18095 12152 18107 12155
rect 18708 12152 18736 12260
rect 20806 12248 20812 12260
rect 20864 12248 20870 12300
rect 22940 12297 22968 12328
rect 23661 12325 23673 12328
rect 23707 12325 23719 12359
rect 23661 12319 23719 12325
rect 22925 12291 22983 12297
rect 22925 12257 22937 12291
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 23014 12248 23020 12300
rect 23072 12248 23078 12300
rect 23109 12291 23167 12297
rect 23109 12257 23121 12291
rect 23155 12288 23167 12291
rect 23290 12288 23296 12300
rect 23155 12260 23296 12288
rect 23155 12257 23167 12260
rect 23109 12251 23167 12257
rect 18966 12180 18972 12232
rect 19024 12180 19030 12232
rect 19334 12180 19340 12232
rect 19392 12180 19398 12232
rect 23124 12220 23152 12251
rect 23290 12248 23296 12260
rect 23348 12288 23354 12300
rect 23768 12297 23796 12396
rect 24302 12384 24308 12436
rect 24360 12424 24366 12436
rect 25130 12424 25136 12436
rect 24360 12396 25136 12424
rect 24360 12384 24366 12396
rect 25130 12384 25136 12396
rect 25188 12384 25194 12436
rect 25222 12384 25228 12436
rect 25280 12384 25286 12436
rect 26326 12384 26332 12436
rect 26384 12424 26390 12436
rect 26602 12424 26608 12436
rect 26384 12396 26608 12424
rect 26384 12384 26390 12396
rect 26602 12384 26608 12396
rect 26660 12384 26666 12436
rect 26786 12384 26792 12436
rect 26844 12424 26850 12436
rect 26881 12427 26939 12433
rect 26881 12424 26893 12427
rect 26844 12396 26893 12424
rect 26844 12384 26850 12396
rect 26881 12393 26893 12396
rect 26927 12393 26939 12427
rect 26881 12387 26939 12393
rect 29549 12427 29607 12433
rect 29549 12393 29561 12427
rect 29595 12424 29607 12427
rect 29730 12424 29736 12436
rect 29595 12396 29736 12424
rect 29595 12393 29607 12396
rect 29549 12387 29607 12393
rect 29730 12384 29736 12396
rect 29788 12384 29794 12436
rect 30193 12427 30251 12433
rect 30193 12393 30205 12427
rect 30239 12424 30251 12427
rect 31754 12424 31760 12436
rect 30239 12396 31760 12424
rect 30239 12393 30251 12396
rect 30193 12387 30251 12393
rect 31754 12384 31760 12396
rect 31812 12424 31818 12436
rect 32490 12424 32496 12436
rect 31812 12396 32496 12424
rect 31812 12384 31818 12396
rect 32490 12384 32496 12396
rect 32548 12384 32554 12436
rect 32674 12384 32680 12436
rect 32732 12424 32738 12436
rect 32950 12424 32956 12436
rect 32732 12396 32956 12424
rect 32732 12384 32738 12396
rect 32950 12384 32956 12396
rect 33008 12384 33014 12436
rect 24412 12328 28994 12356
rect 23569 12291 23627 12297
rect 23569 12288 23581 12291
rect 23348 12260 23581 12288
rect 23348 12248 23354 12260
rect 23569 12257 23581 12260
rect 23615 12257 23627 12291
rect 23569 12251 23627 12257
rect 23753 12291 23811 12297
rect 23753 12257 23765 12291
rect 23799 12257 23811 12291
rect 23753 12251 23811 12257
rect 24412 12232 24440 12328
rect 24762 12248 24768 12300
rect 24820 12288 24826 12300
rect 25777 12291 25835 12297
rect 25777 12288 25789 12291
rect 24820 12260 25789 12288
rect 24820 12248 24826 12260
rect 25777 12257 25789 12260
rect 25823 12257 25835 12291
rect 25777 12251 25835 12257
rect 26234 12248 26240 12300
rect 26292 12248 26298 12300
rect 26326 12248 26332 12300
rect 26384 12288 26390 12300
rect 27798 12288 27804 12300
rect 26384 12260 27804 12288
rect 26384 12248 26390 12260
rect 27798 12248 27804 12260
rect 27856 12248 27862 12300
rect 28966 12288 28994 12328
rect 30285 12291 30343 12297
rect 30285 12288 30297 12291
rect 28966 12260 30297 12288
rect 30285 12257 30297 12260
rect 30331 12288 30343 12291
rect 30331 12260 30512 12288
rect 30331 12257 30343 12260
rect 30285 12251 30343 12257
rect 30484 12232 30512 12260
rect 32306 12248 32312 12300
rect 32364 12288 32370 12300
rect 32364 12260 33272 12288
rect 32364 12248 32370 12260
rect 33244 12232 33272 12260
rect 21560 12192 23152 12220
rect 18095 12124 18736 12152
rect 18877 12155 18935 12161
rect 18095 12121 18107 12124
rect 18049 12115 18107 12121
rect 18877 12121 18889 12155
rect 18923 12152 18935 12155
rect 20070 12152 20076 12164
rect 18923 12124 20076 12152
rect 18923 12121 18935 12124
rect 18877 12115 18935 12121
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 21450 12112 21456 12164
rect 21508 12152 21514 12164
rect 21560 12161 21588 12192
rect 23198 12180 23204 12232
rect 23256 12180 23262 12232
rect 23477 12223 23535 12229
rect 23477 12220 23489 12223
rect 23308 12192 23489 12220
rect 21818 12161 21824 12164
rect 21545 12155 21603 12161
rect 21545 12152 21557 12155
rect 21508 12124 21557 12152
rect 21508 12112 21514 12124
rect 21545 12121 21557 12124
rect 21591 12121 21603 12155
rect 21545 12115 21603 12121
rect 21761 12155 21824 12161
rect 21761 12121 21773 12155
rect 21807 12121 21824 12155
rect 21761 12115 21824 12121
rect 21818 12112 21824 12115
rect 21876 12112 21882 12164
rect 23014 12112 23020 12164
rect 23072 12152 23078 12164
rect 23308 12152 23336 12192
rect 23477 12189 23489 12192
rect 23523 12189 23535 12223
rect 23477 12183 23535 12189
rect 23842 12180 23848 12232
rect 23900 12220 23906 12232
rect 24394 12220 24400 12232
rect 23900 12192 24400 12220
rect 23900 12180 23906 12192
rect 24394 12180 24400 12192
rect 24452 12180 24458 12232
rect 25593 12223 25651 12229
rect 25593 12189 25605 12223
rect 25639 12220 25651 12223
rect 26418 12220 26424 12232
rect 25639 12192 26424 12220
rect 25639 12189 25651 12192
rect 25593 12183 25651 12189
rect 26418 12180 26424 12192
rect 26476 12180 26482 12232
rect 27154 12180 27160 12232
rect 27212 12220 27218 12232
rect 29825 12223 29883 12229
rect 29825 12220 29837 12223
rect 27212 12192 29837 12220
rect 27212 12180 27218 12192
rect 29825 12189 29837 12192
rect 29871 12189 29883 12223
rect 29825 12183 29883 12189
rect 30006 12180 30012 12232
rect 30064 12180 30070 12232
rect 30377 12223 30435 12229
rect 30377 12220 30389 12223
rect 30116 12192 30389 12220
rect 29917 12155 29975 12161
rect 29917 12152 29929 12155
rect 23072 12124 23336 12152
rect 23400 12124 29929 12152
rect 23072 12112 23078 12124
rect 17589 12087 17647 12093
rect 17589 12053 17601 12087
rect 17635 12053 17647 12087
rect 17589 12047 17647 12053
rect 17678 12044 17684 12096
rect 17736 12084 17742 12096
rect 17957 12087 18015 12093
rect 17957 12084 17969 12087
rect 17736 12056 17969 12084
rect 17736 12044 17742 12056
rect 17957 12053 17969 12056
rect 18003 12053 18015 12087
rect 17957 12047 18015 12053
rect 19426 12044 19432 12096
rect 19484 12084 19490 12096
rect 19521 12087 19579 12093
rect 19521 12084 19533 12087
rect 19484 12056 19533 12084
rect 19484 12044 19490 12056
rect 19521 12053 19533 12056
rect 19567 12053 19579 12087
rect 19521 12047 19579 12053
rect 21913 12087 21971 12093
rect 21913 12053 21925 12087
rect 21959 12084 21971 12087
rect 22370 12084 22376 12096
rect 21959 12056 22376 12084
rect 21959 12053 21971 12056
rect 21913 12047 21971 12053
rect 22370 12044 22376 12056
rect 22428 12044 22434 12096
rect 23400 12093 23428 12124
rect 29917 12121 29929 12124
rect 29963 12121 29975 12155
rect 29917 12115 29975 12121
rect 23385 12087 23443 12093
rect 23385 12053 23397 12087
rect 23431 12053 23443 12087
rect 23385 12047 23443 12053
rect 25685 12087 25743 12093
rect 25685 12053 25697 12087
rect 25731 12084 25743 12087
rect 25774 12084 25780 12096
rect 25731 12056 25780 12084
rect 25731 12053 25743 12056
rect 25685 12047 25743 12053
rect 25774 12044 25780 12056
rect 25832 12084 25838 12096
rect 26513 12087 26571 12093
rect 26513 12084 26525 12087
rect 25832 12056 26525 12084
rect 25832 12044 25838 12056
rect 26513 12053 26525 12056
rect 26559 12053 26571 12087
rect 26513 12047 26571 12053
rect 26602 12044 26608 12096
rect 26660 12084 26666 12096
rect 28442 12084 28448 12096
rect 26660 12056 28448 12084
rect 26660 12044 26666 12056
rect 28442 12044 28448 12056
rect 28500 12044 28506 12096
rect 28810 12044 28816 12096
rect 28868 12084 28874 12096
rect 30116 12084 30144 12192
rect 30377 12189 30389 12192
rect 30423 12189 30435 12223
rect 30377 12183 30435 12189
rect 30466 12180 30472 12232
rect 30524 12180 30530 12232
rect 30561 12223 30619 12229
rect 30561 12189 30573 12223
rect 30607 12189 30619 12223
rect 30561 12183 30619 12189
rect 30576 12152 30604 12183
rect 33042 12180 33048 12232
rect 33100 12220 33106 12232
rect 33137 12223 33195 12229
rect 33137 12220 33149 12223
rect 33100 12192 33149 12220
rect 33100 12180 33106 12192
rect 33137 12189 33149 12192
rect 33183 12189 33195 12223
rect 33137 12183 33195 12189
rect 33226 12180 33232 12232
rect 33284 12220 33290 12232
rect 33505 12223 33563 12229
rect 33505 12220 33517 12223
rect 33284 12192 33517 12220
rect 33284 12180 33290 12192
rect 33505 12189 33517 12192
rect 33551 12189 33563 12223
rect 33505 12183 33563 12189
rect 30392 12124 30604 12152
rect 30392 12096 30420 12124
rect 28868 12056 30144 12084
rect 28868 12044 28874 12056
rect 30374 12044 30380 12096
rect 30432 12044 30438 12096
rect 30466 12044 30472 12096
rect 30524 12044 30530 12096
rect 32582 12044 32588 12096
rect 32640 12084 32646 12096
rect 33137 12087 33195 12093
rect 33137 12084 33149 12087
rect 32640 12056 33149 12084
rect 32640 12044 32646 12056
rect 33137 12053 33149 12056
rect 33183 12053 33195 12087
rect 33137 12047 33195 12053
rect 1104 11994 38272 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38272 11994
rect 1104 11920 38272 11942
rect 8754 11840 8760 11892
rect 8812 11880 8818 11892
rect 9306 11880 9312 11892
rect 8812 11852 9312 11880
rect 8812 11840 8818 11852
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 12250 11880 12256 11892
rect 11388 11852 12256 11880
rect 11388 11840 11394 11852
rect 12250 11840 12256 11852
rect 12308 11880 12314 11892
rect 12308 11852 12940 11880
rect 12308 11840 12314 11852
rect 12529 11815 12587 11821
rect 12529 11812 12541 11815
rect 11808 11784 12541 11812
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1489 11747 1547 11753
rect 1489 11744 1501 11747
rect 992 11716 1501 11744
rect 992 11704 998 11716
rect 1489 11713 1501 11716
rect 1535 11713 1547 11747
rect 1489 11707 1547 11713
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 8202 11744 8208 11756
rect 1719 11716 8208 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 10686 11744 10692 11756
rect 9364 11716 10692 11744
rect 9364 11704 9370 11716
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 10778 11704 10784 11756
rect 10836 11704 10842 11756
rect 10318 11636 10324 11688
rect 10376 11676 10382 11688
rect 10870 11676 10876 11688
rect 10376 11648 10876 11676
rect 10376 11636 10382 11648
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 9582 11568 9588 11620
rect 9640 11608 9646 11620
rect 11808 11608 11836 11784
rect 12529 11781 12541 11784
rect 12575 11781 12587 11815
rect 12912 11812 12940 11852
rect 14458 11840 14464 11892
rect 14516 11880 14522 11892
rect 21266 11880 21272 11892
rect 14516 11852 21272 11880
rect 14516 11840 14522 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 22186 11840 22192 11892
rect 22244 11880 22250 11892
rect 22646 11880 22652 11892
rect 22244 11852 22652 11880
rect 22244 11840 22250 11852
rect 22646 11840 22652 11852
rect 22704 11840 22710 11892
rect 24390 11883 24448 11889
rect 24390 11849 24402 11883
rect 24436 11880 24448 11883
rect 27154 11880 27160 11892
rect 24436 11852 27160 11880
rect 24436 11849 24448 11852
rect 24390 11843 24448 11849
rect 27154 11840 27160 11852
rect 27212 11840 27218 11892
rect 27614 11840 27620 11892
rect 27672 11840 27678 11892
rect 29086 11840 29092 11892
rect 29144 11880 29150 11892
rect 29273 11883 29331 11889
rect 29273 11880 29285 11883
rect 29144 11852 29285 11880
rect 29144 11840 29150 11852
rect 29273 11849 29285 11852
rect 29319 11849 29331 11883
rect 29273 11843 29331 11849
rect 29362 11840 29368 11892
rect 29420 11840 29426 11892
rect 29733 11883 29791 11889
rect 29733 11849 29745 11883
rect 29779 11880 29791 11883
rect 30374 11880 30380 11892
rect 29779 11852 30380 11880
rect 29779 11849 29791 11852
rect 29733 11843 29791 11849
rect 30374 11840 30380 11852
rect 30432 11840 30438 11892
rect 32401 11883 32459 11889
rect 32401 11849 32413 11883
rect 32447 11880 32459 11883
rect 32674 11880 32680 11892
rect 32447 11852 32680 11880
rect 32447 11849 32459 11852
rect 32401 11843 32459 11849
rect 32674 11840 32680 11852
rect 32732 11840 32738 11892
rect 12912 11784 13018 11812
rect 12529 11775 12587 11781
rect 15654 11772 15660 11824
rect 15712 11812 15718 11824
rect 15712 11784 16160 11812
rect 15712 11772 15718 11784
rect 11882 11704 11888 11756
rect 11940 11704 11946 11756
rect 11974 11704 11980 11756
rect 12032 11704 12038 11756
rect 14826 11704 14832 11756
rect 14884 11744 14890 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 14884 11716 15945 11744
rect 14884 11704 14890 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 11900 11676 11928 11704
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 11900 11648 12265 11676
rect 12253 11645 12265 11648
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 12894 11636 12900 11688
rect 12952 11676 12958 11688
rect 14274 11676 14280 11688
rect 12952 11648 14280 11676
rect 12952 11636 12958 11648
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 12161 11611 12219 11617
rect 12161 11608 12173 11611
rect 9640 11580 10456 11608
rect 11808 11580 12173 11608
rect 9640 11568 9646 11580
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 8294 11540 8300 11552
rect 3660 11512 8300 11540
rect 3660 11500 3666 11512
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 10318 11500 10324 11552
rect 10376 11500 10382 11552
rect 10428 11540 10456 11580
rect 12161 11577 12173 11580
rect 12207 11577 12219 11611
rect 12161 11571 12219 11577
rect 14844 11540 14872 11704
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15562 11676 15568 11688
rect 15344 11648 15568 11676
rect 15344 11636 15350 11648
rect 15562 11636 15568 11648
rect 15620 11636 15626 11688
rect 16132 11685 16160 11784
rect 18874 11772 18880 11824
rect 18932 11772 18938 11824
rect 21818 11772 21824 11824
rect 21876 11812 21882 11824
rect 22278 11812 22284 11824
rect 21876 11784 22284 11812
rect 21876 11772 21882 11784
rect 22278 11772 22284 11784
rect 22336 11772 22342 11824
rect 26602 11812 26608 11824
rect 23584 11784 24900 11812
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 17604 11716 18613 11744
rect 16025 11679 16083 11685
rect 16025 11645 16037 11679
rect 16071 11645 16083 11679
rect 16025 11639 16083 11645
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11645 16175 11679
rect 16117 11639 16175 11645
rect 16040 11608 16068 11639
rect 17604 11620 17632 11716
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 18785 11747 18843 11753
rect 18785 11713 18797 11747
rect 18831 11744 18843 11747
rect 18892 11744 18920 11772
rect 23584 11756 23612 11784
rect 18831 11716 18920 11744
rect 18831 11713 18843 11716
rect 18785 11707 18843 11713
rect 23566 11704 23572 11756
rect 23624 11704 23630 11756
rect 23753 11747 23811 11753
rect 23753 11713 23765 11747
rect 23799 11744 23811 11747
rect 24118 11744 24124 11756
rect 23799 11716 24124 11744
rect 23799 11713 23811 11716
rect 23753 11707 23811 11713
rect 24118 11704 24124 11716
rect 24176 11704 24182 11756
rect 24210 11704 24216 11756
rect 24268 11704 24274 11756
rect 24305 11747 24363 11753
rect 24305 11713 24317 11747
rect 24351 11744 24363 11747
rect 24394 11744 24400 11756
rect 24351 11716 24400 11744
rect 24351 11713 24363 11716
rect 24305 11707 24363 11713
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 24581 11747 24639 11753
rect 24581 11713 24593 11747
rect 24627 11744 24639 11747
rect 24670 11744 24676 11756
rect 24627 11716 24676 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 23474 11636 23480 11688
rect 23532 11676 23538 11688
rect 23934 11676 23940 11688
rect 23532 11648 23940 11676
rect 23532 11636 23538 11648
rect 23934 11636 23940 11648
rect 23992 11636 23998 11688
rect 17586 11608 17592 11620
rect 16040 11580 17592 11608
rect 17586 11568 17592 11580
rect 17644 11568 17650 11620
rect 18690 11568 18696 11620
rect 18748 11568 18754 11620
rect 22094 11568 22100 11620
rect 22152 11608 22158 11620
rect 24504 11608 24532 11707
rect 24670 11704 24676 11716
rect 24728 11704 24734 11756
rect 24762 11704 24768 11756
rect 24820 11704 24826 11756
rect 24872 11753 24900 11784
rect 25056 11784 26608 11812
rect 25056 11756 25084 11784
rect 26602 11772 26608 11784
rect 26660 11772 26666 11824
rect 27430 11812 27436 11824
rect 27080 11784 27436 11812
rect 24857 11747 24915 11753
rect 24857 11713 24869 11747
rect 24903 11713 24915 11747
rect 24857 11707 24915 11713
rect 25038 11704 25044 11756
rect 25096 11704 25102 11756
rect 24949 11679 25007 11685
rect 24949 11645 24961 11679
rect 24995 11676 25007 11679
rect 26418 11676 26424 11688
rect 24995 11648 26424 11676
rect 24995 11645 25007 11648
rect 24949 11639 25007 11645
rect 26418 11636 26424 11648
rect 26476 11636 26482 11688
rect 24581 11611 24639 11617
rect 24581 11608 24593 11611
rect 22152 11580 24593 11608
rect 22152 11568 22158 11580
rect 24581 11577 24593 11580
rect 24627 11577 24639 11611
rect 27080 11608 27108 11784
rect 27430 11772 27436 11784
rect 27488 11772 27494 11824
rect 27632 11812 27660 11840
rect 27632 11784 27736 11812
rect 27663 11781 27736 11784
rect 27430 11769 27488 11772
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 27172 11676 27200 11707
rect 27338 11704 27344 11756
rect 27396 11704 27402 11756
rect 27430 11735 27442 11769
rect 27476 11735 27488 11769
rect 27663 11747 27675 11781
rect 27709 11750 27736 11781
rect 27798 11772 27804 11824
rect 27856 11812 27862 11824
rect 27893 11815 27951 11821
rect 27893 11812 27905 11815
rect 27856 11784 27905 11812
rect 27856 11772 27862 11784
rect 27893 11781 27905 11784
rect 27939 11812 27951 11815
rect 27982 11812 27988 11824
rect 27939 11784 27988 11812
rect 27939 11781 27951 11784
rect 27893 11775 27951 11781
rect 27982 11772 27988 11784
rect 28040 11772 28046 11824
rect 29380 11812 29408 11840
rect 30193 11815 30251 11821
rect 30193 11812 30205 11815
rect 29380 11784 30205 11812
rect 30193 11781 30205 11784
rect 30239 11781 30251 11815
rect 32214 11812 32220 11824
rect 30193 11775 30251 11781
rect 30300 11784 32220 11812
rect 30300 11756 30328 11784
rect 32214 11772 32220 11784
rect 32272 11812 32278 11824
rect 32272 11784 32720 11812
rect 32272 11772 32278 11784
rect 27709 11747 27721 11750
rect 27663 11741 27721 11747
rect 27430 11729 27488 11735
rect 28810 11704 28816 11756
rect 28868 11704 28874 11756
rect 28994 11704 29000 11756
rect 29052 11744 29058 11756
rect 29457 11747 29515 11753
rect 29457 11744 29469 11747
rect 29052 11716 29469 11744
rect 29052 11704 29058 11716
rect 29457 11713 29469 11716
rect 29503 11713 29515 11747
rect 29457 11707 29515 11713
rect 29730 11704 29736 11756
rect 29788 11744 29794 11756
rect 29917 11747 29975 11753
rect 29917 11744 29929 11747
rect 29788 11716 29929 11744
rect 29788 11704 29794 11716
rect 29917 11713 29929 11716
rect 29963 11713 29975 11747
rect 29917 11707 29975 11713
rect 30282 11704 30288 11756
rect 30340 11704 30346 11756
rect 30466 11704 30472 11756
rect 30524 11744 30530 11756
rect 30561 11747 30619 11753
rect 30561 11744 30573 11747
rect 30524 11716 30573 11744
rect 30524 11704 30530 11716
rect 30561 11713 30573 11716
rect 30607 11713 30619 11747
rect 30561 11707 30619 11713
rect 32582 11704 32588 11756
rect 32640 11704 32646 11756
rect 32692 11753 32720 11784
rect 32677 11747 32735 11753
rect 32677 11713 32689 11747
rect 32723 11744 32735 11747
rect 33686 11744 33692 11756
rect 32723 11716 33692 11744
rect 32723 11713 32735 11716
rect 32677 11707 32735 11713
rect 33686 11704 33692 11716
rect 33744 11704 33750 11756
rect 28828 11676 28856 11704
rect 29549 11679 29607 11685
rect 29549 11676 29561 11679
rect 27172 11648 27568 11676
rect 28828 11648 29561 11676
rect 27540 11620 27568 11648
rect 29549 11645 29561 11648
rect 29595 11645 29607 11679
rect 29549 11639 29607 11645
rect 29822 11636 29828 11688
rect 29880 11636 29886 11688
rect 30650 11636 30656 11688
rect 30708 11636 30714 11688
rect 27154 11608 27160 11620
rect 27080 11580 27160 11608
rect 24581 11571 24639 11577
rect 27154 11568 27160 11580
rect 27212 11568 27218 11620
rect 27522 11568 27528 11620
rect 27580 11568 27586 11620
rect 27890 11568 27896 11620
rect 27948 11608 27954 11620
rect 34606 11608 34612 11620
rect 27948 11580 34612 11608
rect 27948 11568 27954 11580
rect 34606 11568 34612 11580
rect 34664 11568 34670 11620
rect 10428 11512 14872 11540
rect 15562 11500 15568 11552
rect 15620 11500 15626 11552
rect 19242 11500 19248 11552
rect 19300 11540 19306 11552
rect 23474 11540 23480 11552
rect 19300 11512 23480 11540
rect 19300 11500 19306 11512
rect 23474 11500 23480 11512
rect 23532 11500 23538 11552
rect 23569 11543 23627 11549
rect 23569 11509 23581 11543
rect 23615 11540 23627 11543
rect 25774 11540 25780 11552
rect 23615 11512 25780 11540
rect 23615 11509 23627 11512
rect 23569 11503 23627 11509
rect 25774 11500 25780 11512
rect 25832 11500 25838 11552
rect 26878 11500 26884 11552
rect 26936 11540 26942 11552
rect 26973 11543 27031 11549
rect 26973 11540 26985 11543
rect 26936 11512 26985 11540
rect 26936 11500 26942 11512
rect 26973 11509 26985 11512
rect 27019 11540 27031 11543
rect 27430 11540 27436 11552
rect 27019 11512 27436 11540
rect 27019 11509 27031 11512
rect 26973 11503 27031 11509
rect 27430 11500 27436 11512
rect 27488 11500 27494 11552
rect 27706 11500 27712 11552
rect 27764 11500 27770 11552
rect 27982 11500 27988 11552
rect 28040 11540 28046 11552
rect 30282 11540 30288 11552
rect 28040 11512 30288 11540
rect 28040 11500 28046 11512
rect 30282 11500 30288 11512
rect 30340 11500 30346 11552
rect 30374 11500 30380 11552
rect 30432 11540 30438 11552
rect 30837 11543 30895 11549
rect 30837 11540 30849 11543
rect 30432 11512 30849 11540
rect 30432 11500 30438 11512
rect 30837 11509 30849 11512
rect 30883 11509 30895 11543
rect 30837 11503 30895 11509
rect 1104 11450 38272 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38272 11450
rect 1104 11376 38272 11398
rect 3142 11296 3148 11348
rect 3200 11296 3206 11348
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 5718 11336 5724 11348
rect 3476 11308 5724 11336
rect 3476 11296 3482 11308
rect 5718 11296 5724 11308
rect 5776 11296 5782 11348
rect 7834 11296 7840 11348
rect 7892 11296 7898 11348
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 9122 11336 9128 11348
rect 8536 11308 9128 11336
rect 8536 11296 8542 11308
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 10318 11336 10324 11348
rect 9784 11308 10324 11336
rect 3878 11228 3884 11280
rect 3936 11268 3942 11280
rect 3936 11240 4384 11268
rect 3936 11228 3942 11240
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 4062 11200 4068 11212
rect 1443 11172 4068 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4356 11209 4384 11240
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11200 4399 11203
rect 5626 11200 5632 11212
rect 4387 11172 5632 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 7852 11200 7880 11296
rect 8021 11271 8079 11277
rect 8021 11237 8033 11271
rect 8067 11237 8079 11271
rect 8846 11268 8852 11280
rect 8021 11231 8079 11237
rect 8312 11240 8852 11268
rect 7668 11172 7880 11200
rect 5902 11092 5908 11144
rect 5960 11092 5966 11144
rect 6086 11092 6092 11144
rect 6144 11092 6150 11144
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 1670 11024 1676 11076
rect 1728 11024 1734 11076
rect 2958 11064 2964 11076
rect 2898 11036 2964 11064
rect 2958 11024 2964 11036
rect 3016 11064 3022 11076
rect 3878 11064 3884 11076
rect 3016 11036 3884 11064
rect 3016 11024 3022 11036
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 4157 11067 4215 11073
rect 4157 11033 4169 11067
rect 4203 11064 4215 11067
rect 5810 11064 5816 11076
rect 4203 11036 5816 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 7392 11064 7420 11095
rect 7466 11092 7472 11144
rect 7524 11092 7530 11144
rect 7668 11141 7696 11172
rect 7653 11135 7711 11141
rect 7653 11101 7665 11135
rect 7699 11101 7711 11135
rect 7653 11095 7711 11101
rect 7745 11135 7803 11141
rect 7745 11101 7757 11135
rect 7791 11132 7803 11135
rect 8036 11132 8064 11231
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 8312 11209 8340 11240
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 9306 11228 9312 11280
rect 9364 11228 9370 11280
rect 9582 11228 9588 11280
rect 9640 11228 9646 11280
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 8260 11172 8309 11200
rect 8260 11160 8266 11172
rect 8297 11169 8309 11172
rect 8343 11169 8355 11203
rect 9217 11203 9275 11209
rect 9217 11200 9229 11203
rect 8297 11163 8355 11169
rect 9048 11172 9229 11200
rect 7791 11104 8064 11132
rect 7791 11101 7803 11104
rect 7745 11095 7803 11101
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 9048 11132 9076 11172
rect 9217 11169 9229 11172
rect 9263 11200 9275 11203
rect 9600 11200 9628 11228
rect 9263 11172 9628 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 8628 11104 9076 11132
rect 8628 11092 8634 11104
rect 9122 11092 9128 11144
rect 9180 11092 9186 11144
rect 9398 11092 9404 11144
rect 9456 11092 9462 11144
rect 9784 11141 9812 11308
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 12437 11339 12495 11345
rect 12437 11336 12449 11339
rect 12032 11308 12449 11336
rect 12032 11296 12038 11308
rect 12437 11305 12449 11308
rect 12483 11305 12495 11339
rect 14458 11336 14464 11348
rect 12437 11299 12495 11305
rect 12820 11308 14464 11336
rect 9953 11271 10011 11277
rect 9953 11237 9965 11271
rect 9999 11268 10011 11271
rect 12820 11268 12848 11308
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 17586 11296 17592 11348
rect 17644 11296 17650 11348
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 23474 11336 23480 11348
rect 19484 11308 23480 11336
rect 19484 11296 19490 11308
rect 23474 11296 23480 11308
rect 23532 11296 23538 11348
rect 25038 11296 25044 11348
rect 25096 11296 25102 11348
rect 28905 11339 28963 11345
rect 28905 11305 28917 11339
rect 28951 11336 28963 11339
rect 29178 11336 29184 11348
rect 28951 11308 29184 11336
rect 28951 11305 28963 11308
rect 28905 11299 28963 11305
rect 29178 11296 29184 11308
rect 29236 11296 29242 11348
rect 29273 11339 29331 11345
rect 29273 11305 29285 11339
rect 29319 11336 29331 11339
rect 30098 11336 30104 11348
rect 29319 11308 30104 11336
rect 29319 11305 29331 11308
rect 29273 11299 29331 11305
rect 30098 11296 30104 11308
rect 30156 11296 30162 11348
rect 30374 11296 30380 11348
rect 30432 11296 30438 11348
rect 30650 11296 30656 11348
rect 30708 11336 30714 11348
rect 31389 11339 31447 11345
rect 31389 11336 31401 11339
rect 30708 11308 31401 11336
rect 30708 11296 30714 11308
rect 31389 11305 31401 11308
rect 31435 11305 31447 11339
rect 31389 11299 31447 11305
rect 32122 11296 32128 11348
rect 32180 11296 32186 11348
rect 32674 11296 32680 11348
rect 32732 11296 32738 11348
rect 34606 11296 34612 11348
rect 34664 11296 34670 11348
rect 9999 11240 10180 11268
rect 9999 11237 10011 11240
rect 9953 11231 10011 11237
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9916 11172 10057 11200
rect 9916 11160 9922 11172
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10152 11200 10180 11240
rect 12406 11240 12848 11268
rect 14093 11271 14151 11277
rect 10321 11203 10379 11209
rect 10321 11200 10333 11203
rect 10152 11172 10333 11200
rect 10045 11163 10103 11169
rect 10321 11169 10333 11172
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 10778 11160 10784 11212
rect 10836 11200 10842 11212
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 10836 11172 11805 11200
rect 10836 11160 10842 11172
rect 11793 11169 11805 11172
rect 11839 11200 11851 11203
rect 12406 11200 12434 11240
rect 14093 11237 14105 11271
rect 14139 11237 14151 11271
rect 15286 11268 15292 11280
rect 14093 11231 14151 11237
rect 14752 11240 15292 11268
rect 11839 11172 12434 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 12894 11160 12900 11212
rect 12952 11160 12958 11212
rect 13081 11203 13139 11209
rect 13081 11169 13093 11203
rect 13127 11200 13139 11203
rect 13127 11172 13492 11200
rect 13127 11169 13139 11172
rect 13081 11163 13139 11169
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 13096 11132 13124 11163
rect 12676 11104 13124 11132
rect 12676 11092 12682 11104
rect 7558 11064 7564 11076
rect 7392 11036 7564 11064
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 7834 11024 7840 11076
rect 7892 11064 7898 11076
rect 7929 11067 7987 11073
rect 7929 11064 7941 11067
rect 7892 11036 7941 11064
rect 7892 11024 7898 11036
rect 7929 11033 7941 11036
rect 7975 11033 7987 11067
rect 7929 11027 7987 11033
rect 8110 11024 8116 11076
rect 8168 11064 8174 11076
rect 8941 11067 8999 11073
rect 8941 11064 8953 11067
rect 8168 11036 8953 11064
rect 8168 11024 8174 11036
rect 8941 11033 8953 11036
rect 8987 11033 8999 11067
rect 8941 11027 8999 11033
rect 11330 11024 11336 11076
rect 11388 11024 11394 11076
rect 12802 11024 12808 11076
rect 12860 11064 12866 11076
rect 13354 11064 13360 11076
rect 12860 11036 13360 11064
rect 12860 11024 12866 11036
rect 13354 11024 13360 11036
rect 13412 11024 13418 11076
rect 13464 11064 13492 11172
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 14108 11132 14136 11231
rect 14752 11209 14780 11240
rect 15286 11228 15292 11240
rect 15344 11228 15350 11280
rect 15749 11271 15807 11277
rect 15749 11237 15761 11271
rect 15795 11268 15807 11271
rect 15795 11240 15976 11268
rect 15795 11237 15807 11240
rect 15749 11231 15807 11237
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 13771 11104 14136 11132
rect 14200 11172 14749 11200
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 14200 11064 14228 11172
rect 14737 11169 14749 11172
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 14826 11160 14832 11212
rect 14884 11160 14890 11212
rect 15948 11200 15976 11240
rect 18782 11228 18788 11280
rect 18840 11228 18846 11280
rect 19242 11228 19248 11280
rect 19300 11228 19306 11280
rect 16117 11203 16175 11209
rect 16117 11200 16129 11203
rect 15948 11172 16129 11200
rect 16117 11169 16129 11172
rect 16163 11169 16175 11203
rect 18800 11200 18828 11228
rect 16117 11163 16175 11169
rect 18708 11172 18828 11200
rect 19260 11200 19288 11228
rect 19260 11172 19380 11200
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11132 14519 11135
rect 14844 11132 14872 11160
rect 14507 11104 14872 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 15562 11092 15568 11144
rect 15620 11092 15626 11144
rect 15746 11092 15752 11144
rect 15804 11132 15810 11144
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 15804 11104 15853 11132
rect 15804 11092 15810 11104
rect 15841 11101 15853 11104
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 18601 11135 18659 11141
rect 18601 11132 18613 11135
rect 18288 11104 18613 11132
rect 18288 11092 18294 11104
rect 18601 11101 18613 11104
rect 18647 11101 18659 11135
rect 18601 11095 18659 11101
rect 18417 11067 18475 11073
rect 13464 11036 14228 11064
rect 16500 11036 16606 11064
rect 16500 11008 16528 11036
rect 18417 11033 18429 11067
rect 18463 11064 18475 11067
rect 18708 11064 18736 11172
rect 18785 11135 18843 11141
rect 18785 11101 18797 11135
rect 18831 11132 18843 11135
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18831 11104 19257 11132
rect 18831 11101 18843 11104
rect 18785 11095 18843 11101
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 18463 11036 18736 11064
rect 19352 11064 19380 11172
rect 19444 11132 19472 11296
rect 20254 11228 20260 11280
rect 20312 11228 20318 11280
rect 21818 11228 21824 11280
rect 21876 11228 21882 11280
rect 21913 11271 21971 11277
rect 21913 11237 21925 11271
rect 21959 11268 21971 11271
rect 22278 11268 22284 11280
rect 21959 11240 22284 11268
rect 21959 11237 21971 11240
rect 21913 11231 21971 11237
rect 22278 11228 22284 11240
rect 22336 11228 22342 11280
rect 23566 11268 23572 11280
rect 22388 11240 23572 11268
rect 20272 11200 20300 11228
rect 21836 11200 21864 11228
rect 22388 11212 22416 11240
rect 23566 11228 23572 11240
rect 23624 11228 23630 11280
rect 25056 11268 25084 11296
rect 26602 11268 26608 11280
rect 23768 11240 25084 11268
rect 26344 11240 26608 11268
rect 22370 11200 22376 11212
rect 19996 11172 20300 11200
rect 21376 11172 21864 11200
rect 22204 11172 22376 11200
rect 19996 11141 20024 11172
rect 19889 11135 19947 11141
rect 19889 11132 19901 11135
rect 19444 11104 19901 11132
rect 19889 11101 19901 11104
rect 19935 11101 19947 11135
rect 19889 11095 19947 11101
rect 19981 11135 20039 11141
rect 19981 11101 19993 11135
rect 20027 11101 20039 11135
rect 19981 11095 20039 11101
rect 20070 11092 20076 11144
rect 20128 11092 20134 11144
rect 21376 11141 21404 11172
rect 22204 11141 22232 11172
rect 22370 11160 22376 11172
rect 22428 11160 22434 11212
rect 23106 11200 23112 11212
rect 22480 11172 23112 11200
rect 22480 11141 22508 11172
rect 23106 11160 23112 11172
rect 23164 11160 23170 11212
rect 23768 11209 23796 11240
rect 26344 11212 26372 11240
rect 26602 11228 26608 11240
rect 26660 11228 26666 11280
rect 27062 11228 27068 11280
rect 27120 11268 27126 11280
rect 27120 11240 27292 11268
rect 27120 11228 27126 11240
rect 23753 11203 23811 11209
rect 23753 11169 23765 11203
rect 23799 11169 23811 11203
rect 23753 11163 23811 11169
rect 21361 11135 21419 11141
rect 21361 11101 21373 11135
rect 21407 11101 21419 11135
rect 21637 11135 21695 11141
rect 21637 11132 21649 11135
rect 21361 11095 21419 11101
rect 21468 11104 21649 11132
rect 19521 11067 19579 11073
rect 19521 11064 19533 11067
rect 19352 11036 19533 11064
rect 18463 11033 18475 11036
rect 18417 11027 18475 11033
rect 19521 11033 19533 11036
rect 19567 11033 19579 11067
rect 19521 11027 19579 11033
rect 20257 11067 20315 11073
rect 20257 11033 20269 11067
rect 20303 11064 20315 11067
rect 20990 11064 20996 11076
rect 20303 11036 20996 11064
rect 20303 11033 20315 11036
rect 20257 11027 20315 11033
rect 20990 11024 20996 11036
rect 21048 11064 21054 11076
rect 21468 11064 21496 11104
rect 21637 11101 21649 11104
rect 21683 11101 21695 11135
rect 21637 11095 21695 11101
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11132 21787 11135
rect 22005 11135 22063 11141
rect 22005 11132 22017 11135
rect 21775 11104 22017 11132
rect 21775 11101 21787 11104
rect 21729 11095 21787 11101
rect 22005 11101 22017 11104
rect 22051 11101 22063 11135
rect 22005 11095 22063 11101
rect 22189 11135 22247 11141
rect 22189 11101 22201 11135
rect 22235 11101 22247 11135
rect 22189 11095 22247 11101
rect 22465 11135 22523 11141
rect 22465 11101 22477 11135
rect 22511 11101 22523 11135
rect 22465 11095 22523 11101
rect 23569 11135 23627 11141
rect 23569 11101 23581 11135
rect 23615 11132 23627 11135
rect 23658 11132 23664 11144
rect 23615 11104 23664 11132
rect 23615 11101 23627 11104
rect 23569 11095 23627 11101
rect 23658 11092 23664 11104
rect 23716 11092 23722 11144
rect 21048 11036 21496 11064
rect 21545 11067 21603 11073
rect 21048 11024 21054 11036
rect 21545 11033 21557 11067
rect 21591 11033 21603 11067
rect 22094 11064 22100 11076
rect 21545 11027 21603 11033
rect 21744 11036 22100 11064
rect 3786 10956 3792 11008
rect 3844 10956 3850 11008
rect 4246 10956 4252 11008
rect 4304 10956 4310 11008
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 12342 10996 12348 11008
rect 6788 10968 12348 10996
rect 6788 10956 6794 10968
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 13909 10999 13967 11005
rect 13909 10965 13921 10999
rect 13955 10996 13967 10999
rect 14090 10996 14096 11008
rect 13955 10968 14096 10996
rect 13955 10965 13967 10968
rect 13909 10959 13967 10965
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 14553 10999 14611 11005
rect 14553 10965 14565 10999
rect 14599 10996 14611 10999
rect 15930 10996 15936 11008
rect 14599 10968 15936 10996
rect 14599 10965 14611 10968
rect 14553 10959 14611 10965
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 16482 10956 16488 11008
rect 16540 10956 16546 11008
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 21450 10996 21456 11008
rect 17092 10968 21456 10996
rect 17092 10956 17098 10968
rect 21450 10956 21456 10968
rect 21508 10956 21514 11008
rect 21560 10996 21588 11027
rect 21744 10996 21772 11036
rect 22094 11024 22100 11036
rect 22152 11024 22158 11076
rect 22373 11067 22431 11073
rect 22373 11064 22385 11067
rect 22204 11036 22385 11064
rect 21560 10968 21772 10996
rect 21818 10956 21824 11008
rect 21876 10996 21882 11008
rect 22204 10996 22232 11036
rect 22373 11033 22385 11036
rect 22419 11033 22431 11067
rect 22373 11027 22431 11033
rect 23290 11024 23296 11076
rect 23348 11064 23354 11076
rect 23768 11064 23796 11163
rect 24210 11160 24216 11212
rect 24268 11200 24274 11212
rect 24762 11200 24768 11212
rect 24268 11172 24768 11200
rect 24268 11160 24274 11172
rect 24762 11160 24768 11172
rect 24820 11200 24826 11212
rect 26145 11203 26203 11209
rect 24820 11172 25452 11200
rect 24820 11160 24826 11172
rect 25424 11141 25452 11172
rect 26145 11169 26157 11203
rect 26191 11200 26203 11203
rect 26326 11200 26332 11212
rect 26191 11172 26332 11200
rect 26191 11169 26203 11172
rect 26145 11163 26203 11169
rect 26326 11160 26332 11172
rect 26384 11160 26390 11212
rect 27157 11203 27215 11209
rect 27157 11200 27169 11203
rect 26528 11172 27169 11200
rect 26528 11144 26556 11172
rect 27157 11169 27169 11172
rect 27203 11169 27215 11203
rect 27157 11163 27215 11169
rect 25409 11135 25467 11141
rect 25409 11101 25421 11135
rect 25455 11101 25467 11135
rect 25409 11095 25467 11101
rect 25593 11135 25651 11141
rect 25593 11101 25605 11135
rect 25639 11132 25651 11135
rect 26234 11132 26240 11144
rect 25639 11104 26240 11132
rect 25639 11101 25651 11104
rect 25593 11095 25651 11101
rect 26234 11092 26240 11104
rect 26292 11092 26298 11144
rect 26418 11092 26424 11144
rect 26476 11092 26482 11144
rect 26510 11092 26516 11144
rect 26568 11092 26574 11144
rect 26881 11135 26939 11141
rect 26881 11101 26893 11135
rect 26927 11101 26939 11135
rect 26881 11095 26939 11101
rect 23348 11036 23796 11064
rect 25501 11067 25559 11073
rect 23348 11024 23354 11036
rect 25501 11033 25513 11067
rect 25547 11064 25559 11067
rect 26896 11064 26924 11095
rect 27062 11092 27068 11144
rect 27120 11092 27126 11144
rect 27264 11141 27292 11240
rect 27338 11228 27344 11280
rect 27396 11228 27402 11280
rect 27430 11228 27436 11280
rect 27488 11268 27494 11280
rect 30392 11268 30420 11296
rect 27488 11240 29132 11268
rect 27488 11228 27494 11240
rect 27249 11135 27307 11141
rect 27249 11101 27261 11135
rect 27295 11101 27307 11135
rect 27356 11132 27384 11228
rect 27614 11160 27620 11212
rect 27672 11200 27678 11212
rect 27672 11172 28212 11200
rect 27672 11160 27678 11172
rect 27433 11135 27491 11141
rect 27433 11132 27445 11135
rect 27356 11104 27445 11132
rect 27249 11095 27307 11101
rect 27433 11101 27445 11104
rect 27479 11132 27491 11135
rect 27709 11135 27767 11141
rect 27709 11132 27721 11135
rect 27479 11104 27721 11132
rect 27479 11101 27491 11104
rect 27433 11095 27491 11101
rect 27709 11101 27721 11104
rect 27755 11101 27767 11135
rect 27709 11095 27767 11101
rect 27264 11064 27292 11095
rect 27798 11092 27804 11144
rect 27856 11092 27862 11144
rect 27893 11135 27951 11141
rect 27893 11101 27905 11135
rect 27939 11132 27951 11135
rect 27982 11132 27988 11144
rect 27939 11104 27988 11132
rect 27939 11101 27951 11104
rect 27893 11095 27951 11101
rect 27982 11092 27988 11104
rect 28040 11092 28046 11144
rect 28184 11141 28212 11172
rect 29104 11141 29132 11240
rect 30116 11240 30420 11268
rect 30561 11271 30619 11277
rect 30116 11209 30144 11240
rect 30561 11237 30573 11271
rect 30607 11268 30619 11271
rect 31754 11268 31760 11280
rect 30607 11240 31760 11268
rect 30607 11237 30619 11240
rect 30561 11231 30619 11237
rect 31754 11228 31760 11240
rect 31812 11228 31818 11280
rect 32692 11268 32720 11296
rect 31864 11240 33088 11268
rect 30101 11203 30159 11209
rect 30101 11169 30113 11203
rect 30147 11169 30159 11203
rect 30101 11163 30159 11169
rect 30466 11160 30472 11212
rect 30524 11160 30530 11212
rect 31864 11200 31892 11240
rect 31726 11172 31892 11200
rect 32324 11172 32904 11200
rect 28169 11135 28227 11141
rect 28169 11101 28181 11135
rect 28215 11132 28227 11135
rect 28261 11135 28319 11141
rect 28261 11132 28273 11135
rect 28215 11104 28273 11132
rect 28215 11101 28227 11104
rect 28169 11095 28227 11101
rect 28261 11101 28273 11104
rect 28307 11101 28319 11135
rect 28445 11135 28503 11141
rect 28445 11132 28457 11135
rect 28261 11095 28319 11101
rect 28368 11104 28457 11132
rect 25547 11036 26924 11064
rect 27080 11036 27292 11064
rect 27816 11064 27844 11092
rect 28077 11067 28135 11073
rect 28077 11064 28089 11067
rect 27816 11036 28089 11064
rect 25547 11033 25559 11036
rect 25501 11027 25559 11033
rect 27080 11008 27108 11036
rect 28077 11033 28089 11036
rect 28123 11064 28135 11067
rect 28368 11064 28396 11104
rect 28445 11101 28457 11104
rect 28491 11101 28503 11135
rect 28445 11095 28503 11101
rect 29089 11135 29147 11141
rect 29089 11101 29101 11135
rect 29135 11101 29147 11135
rect 29089 11095 29147 11101
rect 29365 11135 29423 11141
rect 29365 11101 29377 11135
rect 29411 11132 29423 11135
rect 29638 11132 29644 11144
rect 29411 11104 29644 11132
rect 29411 11101 29423 11104
rect 29365 11095 29423 11101
rect 29638 11092 29644 11104
rect 29696 11132 29702 11144
rect 30190 11132 30196 11144
rect 29696 11104 30196 11132
rect 29696 11092 29702 11104
rect 30190 11092 30196 11104
rect 30248 11092 30254 11144
rect 30282 11092 30288 11144
rect 30340 11092 30346 11144
rect 30377 11135 30435 11141
rect 30377 11101 30389 11135
rect 30423 11132 30435 11135
rect 30484 11132 30512 11160
rect 30423 11104 30512 11132
rect 31573 11135 31631 11141
rect 30423 11101 30435 11104
rect 30377 11095 30435 11101
rect 31573 11101 31585 11135
rect 31619 11132 31631 11135
rect 31726 11132 31754 11172
rect 32324 11144 32352 11172
rect 31619 11104 31754 11132
rect 31619 11101 31631 11104
rect 31573 11095 31631 11101
rect 31846 11092 31852 11144
rect 31904 11092 31910 11144
rect 32033 11135 32091 11141
rect 32033 11101 32045 11135
rect 32079 11132 32091 11135
rect 32306 11132 32312 11144
rect 32079 11104 32312 11132
rect 32079 11101 32091 11104
rect 32033 11095 32091 11101
rect 32306 11092 32312 11104
rect 32364 11092 32370 11144
rect 32490 11092 32496 11144
rect 32548 11132 32554 11144
rect 32585 11135 32643 11141
rect 32585 11132 32597 11135
rect 32548 11104 32597 11132
rect 32548 11092 32554 11104
rect 32585 11101 32597 11104
rect 32631 11101 32643 11135
rect 32585 11095 32643 11101
rect 32766 11092 32772 11144
rect 32824 11092 32830 11144
rect 32876 11141 32904 11172
rect 33060 11141 33088 11240
rect 32861 11135 32919 11141
rect 32861 11101 32873 11135
rect 32907 11101 32919 11135
rect 32861 11095 32919 11101
rect 33045 11135 33103 11141
rect 33045 11101 33057 11135
rect 33091 11101 33103 11135
rect 34624 11132 34652 11296
rect 37553 11135 37611 11141
rect 37553 11132 37565 11135
rect 34624 11104 37565 11132
rect 33045 11095 33103 11101
rect 37553 11101 37565 11104
rect 37599 11101 37611 11135
rect 37553 11095 37611 11101
rect 28123 11036 28396 11064
rect 28460 11036 31754 11064
rect 28123 11033 28135 11036
rect 28077 11027 28135 11033
rect 21876 10968 22232 10996
rect 21876 10956 21882 10968
rect 23382 10956 23388 11008
rect 23440 10956 23446 11008
rect 25774 10956 25780 11008
rect 25832 10996 25838 11008
rect 26329 10999 26387 11005
rect 26329 10996 26341 10999
rect 25832 10968 26341 10996
rect 25832 10956 25838 10968
rect 26329 10965 26341 10968
rect 26375 10965 26387 10999
rect 26329 10959 26387 10965
rect 26786 10956 26792 11008
rect 26844 10956 26850 11008
rect 27062 10956 27068 11008
rect 27120 10956 27126 11008
rect 27614 10956 27620 11008
rect 27672 10956 27678 11008
rect 28460 11005 28488 11036
rect 28445 10999 28503 11005
rect 28445 10965 28457 10999
rect 28491 10965 28503 10999
rect 28445 10959 28503 10965
rect 30190 10956 30196 11008
rect 30248 10996 30254 11008
rect 30650 10996 30656 11008
rect 30248 10968 30656 10996
rect 30248 10956 30254 10968
rect 30650 10956 30656 10968
rect 30708 10956 30714 11008
rect 31726 10996 31754 11036
rect 37918 11024 37924 11076
rect 37976 11024 37982 11076
rect 32582 10996 32588 11008
rect 31726 10968 32588 10996
rect 32582 10956 32588 10968
rect 32640 10956 32646 11008
rect 32950 10956 32956 11008
rect 33008 10956 33014 11008
rect 1104 10906 38272 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38272 10906
rect 1104 10832 38272 10854
rect 1670 10752 1676 10804
rect 1728 10792 1734 10804
rect 1765 10795 1823 10801
rect 1765 10792 1777 10795
rect 1728 10764 1777 10792
rect 1728 10752 1734 10764
rect 1765 10761 1777 10764
rect 1811 10761 1823 10795
rect 1765 10755 1823 10761
rect 2777 10795 2835 10801
rect 2777 10761 2789 10795
rect 2823 10792 2835 10795
rect 3786 10792 3792 10804
rect 2823 10764 3792 10792
rect 2823 10761 2835 10764
rect 2777 10755 2835 10761
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 5813 10795 5871 10801
rect 3936 10764 4384 10792
rect 3936 10752 3942 10764
rect 4246 10724 4252 10736
rect 3712 10696 4252 10724
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10656 2007 10659
rect 2685 10659 2743 10665
rect 1995 10628 2360 10656
rect 1995 10625 2007 10628
rect 1949 10619 2007 10625
rect 2332 10529 2360 10628
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 3142 10656 3148 10668
rect 2731 10628 3148 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 3142 10616 3148 10628
rect 3200 10656 3206 10668
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 3200 10628 3341 10656
rect 3200 10616 3206 10628
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10557 3019 10591
rect 2961 10551 3019 10557
rect 2317 10523 2375 10529
rect 2317 10489 2329 10523
rect 2363 10489 2375 10523
rect 2317 10483 2375 10489
rect 2976 10452 3004 10551
rect 3418 10548 3424 10600
rect 3476 10548 3482 10600
rect 3712 10597 3740 10696
rect 4246 10684 4252 10696
rect 4304 10684 4310 10736
rect 4356 10724 4384 10764
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 6086 10792 6092 10804
rect 5859 10764 6092 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 6086 10752 6092 10764
rect 6144 10792 6150 10804
rect 6144 10764 7420 10792
rect 6144 10752 6150 10764
rect 4356 10696 4830 10724
rect 5626 10684 5632 10736
rect 5684 10724 5690 10736
rect 7392 10733 7420 10764
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 8665 10795 8723 10801
rect 8665 10792 8677 10795
rect 8536 10764 8677 10792
rect 8536 10752 8542 10764
rect 8665 10761 8677 10764
rect 8711 10761 8723 10795
rect 8665 10755 8723 10761
rect 9033 10795 9091 10801
rect 9033 10761 9045 10795
rect 9079 10792 9091 10795
rect 9398 10792 9404 10804
rect 9079 10764 9404 10792
rect 9079 10761 9091 10764
rect 9033 10755 9091 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 15746 10792 15752 10804
rect 13924 10764 15752 10792
rect 7377 10727 7435 10733
rect 5684 10696 6960 10724
rect 5684 10684 5690 10696
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5776 10628 6009 10656
rect 5776 10616 5782 10628
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6178 10616 6184 10668
rect 6236 10616 6242 10668
rect 6730 10616 6736 10668
rect 6788 10616 6794 10668
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10557 3755 10591
rect 3697 10551 3755 10557
rect 4062 10548 4068 10600
rect 4120 10548 4126 10600
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10588 4399 10591
rect 4706 10588 4712 10600
rect 4387 10560 4712 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 5810 10548 5816 10600
rect 5868 10548 5874 10600
rect 6932 10597 6960 10696
rect 7377 10693 7389 10727
rect 7423 10693 7435 10727
rect 7377 10687 7435 10693
rect 7561 10727 7619 10733
rect 7561 10693 7573 10727
rect 7607 10724 7619 10727
rect 13924 10724 13952 10764
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 19153 10795 19211 10801
rect 19153 10792 19165 10795
rect 18932 10764 19165 10792
rect 18932 10752 18938 10764
rect 19153 10761 19165 10764
rect 19199 10761 19211 10795
rect 21542 10792 21548 10804
rect 19153 10755 19211 10761
rect 20824 10764 21548 10792
rect 7607 10696 12204 10724
rect 7607 10693 7619 10696
rect 7561 10687 7619 10693
rect 7190 10616 7196 10668
rect 7248 10616 7254 10668
rect 7466 10616 7472 10668
rect 7524 10656 7530 10668
rect 8478 10656 8484 10668
rect 7524 10628 8484 10656
rect 7524 10616 7530 10628
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10588 6147 10591
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6135 10560 6837 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10557 6975 10591
rect 8588 10588 8616 10619
rect 8846 10616 8852 10668
rect 8904 10616 8910 10668
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 8588 10560 9137 10588
rect 6917 10551 6975 10557
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9600 10588 9628 10619
rect 10778 10616 10784 10668
rect 10836 10656 10842 10668
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10836 10628 10977 10656
rect 10836 10616 10842 10628
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 10226 10588 10232 10600
rect 9125 10551 9183 10557
rect 9232 10560 9444 10588
rect 9600 10560 10232 10588
rect 5828 10520 5856 10548
rect 9232 10520 9260 10560
rect 5828 10492 9260 10520
rect 3234 10452 3240 10464
rect 2976 10424 3240 10452
rect 3234 10412 3240 10424
rect 3292 10452 3298 10464
rect 5810 10452 5816 10464
rect 3292 10424 5816 10452
rect 3292 10412 3298 10424
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 6362 10412 6368 10464
rect 6420 10412 6426 10464
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 9309 10455 9367 10461
rect 9309 10452 9321 10455
rect 8352 10424 9321 10452
rect 8352 10412 8358 10424
rect 9309 10421 9321 10424
rect 9355 10421 9367 10455
rect 9416 10452 9444 10560
rect 10226 10548 10232 10560
rect 10284 10548 10290 10600
rect 11057 10591 11115 10597
rect 11057 10588 11069 10591
rect 10980 10560 11069 10588
rect 10597 10455 10655 10461
rect 10597 10452 10609 10455
rect 9416 10424 10609 10452
rect 9309 10415 9367 10421
rect 10597 10421 10609 10424
rect 10643 10421 10655 10455
rect 10980 10452 11008 10560
rect 11057 10557 11069 10560
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 11238 10548 11244 10600
rect 11296 10548 11302 10600
rect 12176 10520 12204 10696
rect 12268 10696 13952 10724
rect 12268 10600 12296 10696
rect 13924 10665 13952 10696
rect 14090 10684 14096 10736
rect 14148 10724 14154 10736
rect 14185 10727 14243 10733
rect 14185 10724 14197 10727
rect 14148 10696 14197 10724
rect 14148 10684 14154 10696
rect 14185 10693 14197 10696
rect 14231 10693 14243 10727
rect 14185 10687 14243 10693
rect 15930 10684 15936 10736
rect 15988 10684 15994 10736
rect 20824 10733 20852 10764
rect 21542 10752 21548 10764
rect 21600 10752 21606 10804
rect 24121 10795 24179 10801
rect 24121 10792 24133 10795
rect 22296 10764 24133 10792
rect 20809 10727 20867 10733
rect 20809 10724 20821 10727
rect 20272 10696 20821 10724
rect 13909 10659 13967 10665
rect 13909 10625 13921 10659
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 15286 10616 15292 10668
rect 15344 10656 15350 10668
rect 16482 10656 16488 10668
rect 15344 10628 16488 10656
rect 15344 10616 15350 10628
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10656 16911 10659
rect 16942 10656 16948 10668
rect 16899 10628 16948 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 12250 10548 12256 10600
rect 12308 10548 12314 10600
rect 17052 10588 17080 10619
rect 17126 10616 17132 10668
rect 17184 10616 17190 10668
rect 17221 10659 17279 10665
rect 17221 10625 17233 10659
rect 17267 10656 17279 10659
rect 18141 10659 18199 10665
rect 17267 10628 18092 10656
rect 17267 10625 17279 10628
rect 17221 10619 17279 10625
rect 13372 10560 17080 10588
rect 13372 10520 13400 10560
rect 12176 10492 13400 10520
rect 17494 10480 17500 10532
rect 17552 10480 17558 10532
rect 18064 10520 18092 10628
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 18230 10656 18236 10668
rect 18187 10628 18236 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 18230 10616 18236 10628
rect 18288 10656 18294 10668
rect 18325 10659 18383 10665
rect 18325 10656 18337 10659
rect 18288 10628 18337 10656
rect 18288 10616 18294 10628
rect 18325 10625 18337 10628
rect 18371 10625 18383 10659
rect 18325 10619 18383 10625
rect 18782 10616 18788 10668
rect 18840 10656 18846 10668
rect 20272 10665 20300 10696
rect 20809 10693 20821 10696
rect 20855 10693 20867 10727
rect 20809 10687 20867 10693
rect 20990 10684 20996 10736
rect 21048 10733 21054 10736
rect 21048 10727 21067 10733
rect 21055 10724 21067 10727
rect 22296 10724 22324 10764
rect 24121 10761 24133 10764
rect 24167 10761 24179 10795
rect 24121 10755 24179 10761
rect 24213 10795 24271 10801
rect 24213 10761 24225 10795
rect 24259 10792 24271 10795
rect 24394 10792 24400 10804
rect 24259 10764 24400 10792
rect 24259 10761 24271 10764
rect 24213 10755 24271 10761
rect 21055 10696 21496 10724
rect 21055 10693 21067 10696
rect 21048 10687 21067 10693
rect 21048 10684 21054 10687
rect 21468 10665 21496 10696
rect 22112 10696 22324 10724
rect 22112 10665 22140 10696
rect 22922 10684 22928 10736
rect 22980 10684 22986 10736
rect 23106 10684 23112 10736
rect 23164 10684 23170 10736
rect 23247 10727 23305 10733
rect 23247 10693 23259 10727
rect 23293 10724 23305 10727
rect 23382 10724 23388 10736
rect 23293 10696 23388 10724
rect 23293 10693 23305 10696
rect 23247 10687 23305 10693
rect 23382 10684 23388 10696
rect 23440 10684 23446 10736
rect 22926 10681 22984 10684
rect 18969 10659 19027 10665
rect 18969 10656 18981 10659
rect 18840 10628 18981 10656
rect 18840 10616 18846 10628
rect 18969 10625 18981 10628
rect 19015 10625 19027 10659
rect 18969 10619 19027 10625
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10625 20315 10659
rect 20257 10619 20315 10625
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10625 21511 10659
rect 22097 10659 22155 10665
rect 22097 10656 22109 10659
rect 21453 10619 21511 10625
rect 21560 10628 22109 10656
rect 21174 10548 21180 10600
rect 21232 10588 21238 10600
rect 21269 10591 21327 10597
rect 21269 10588 21281 10591
rect 21232 10560 21281 10588
rect 21232 10548 21238 10560
rect 21269 10557 21281 10560
rect 21315 10588 21327 10591
rect 21560 10588 21588 10628
rect 22097 10625 22109 10628
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 21315 10560 21588 10588
rect 21315 10557 21327 10560
rect 21269 10551 21327 10557
rect 21634 10548 21640 10600
rect 21692 10548 21698 10600
rect 21910 10548 21916 10600
rect 21968 10588 21974 10600
rect 22204 10588 22232 10619
rect 22370 10616 22376 10668
rect 22428 10616 22434 10668
rect 22462 10616 22468 10668
rect 22520 10616 22526 10668
rect 22830 10616 22836 10668
rect 22888 10616 22894 10668
rect 22926 10647 22938 10681
rect 22972 10647 22984 10681
rect 22926 10641 22984 10647
rect 23017 10659 23075 10665
rect 23017 10625 23029 10659
rect 23063 10656 23075 10659
rect 23474 10656 23480 10668
rect 23063 10628 23336 10656
rect 23063 10625 23075 10628
rect 23017 10619 23075 10625
rect 22848 10588 22876 10616
rect 23308 10600 23336 10628
rect 23400 10628 23480 10656
rect 23106 10588 23112 10600
rect 21968 10560 22140 10588
rect 22204 10560 23112 10588
rect 21968 10548 21974 10560
rect 20806 10520 20812 10532
rect 18064 10492 20812 10520
rect 20806 10480 20812 10492
rect 20864 10480 20870 10532
rect 21818 10480 21824 10532
rect 21876 10520 21882 10532
rect 22112 10520 22140 10560
rect 23106 10548 23112 10560
rect 23164 10548 23170 10600
rect 23290 10548 23296 10600
rect 23348 10548 23354 10600
rect 23400 10597 23428 10628
rect 23474 10616 23480 10628
rect 23532 10656 23538 10668
rect 24228 10656 24256 10755
rect 24394 10752 24400 10764
rect 24452 10752 24458 10804
rect 27614 10752 27620 10804
rect 27672 10752 27678 10804
rect 28166 10752 28172 10804
rect 28224 10792 28230 10804
rect 32217 10795 32275 10801
rect 28224 10764 28580 10792
rect 28224 10752 28230 10764
rect 27632 10724 27660 10752
rect 28442 10724 28448 10736
rect 27172 10696 27660 10724
rect 28276 10696 28448 10724
rect 23532 10628 24256 10656
rect 23532 10616 23538 10628
rect 26786 10616 26792 10668
rect 26844 10656 26850 10668
rect 27172 10665 27200 10696
rect 26973 10659 27031 10665
rect 26973 10656 26985 10659
rect 26844 10628 26985 10656
rect 26844 10616 26850 10628
rect 26973 10625 26985 10628
rect 27019 10625 27031 10659
rect 26973 10619 27031 10625
rect 27157 10659 27215 10665
rect 27157 10625 27169 10659
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 27246 10616 27252 10668
rect 27304 10616 27310 10668
rect 27341 10659 27399 10665
rect 27341 10625 27353 10659
rect 27387 10656 27399 10659
rect 27522 10656 27528 10668
rect 27387 10628 27528 10656
rect 27387 10625 27399 10628
rect 27341 10619 27399 10625
rect 27522 10616 27528 10628
rect 27580 10616 27586 10668
rect 28276 10665 28304 10696
rect 28442 10684 28448 10696
rect 28500 10684 28506 10736
rect 28552 10733 28580 10764
rect 32217 10761 32229 10795
rect 32263 10792 32275 10795
rect 32306 10792 32312 10804
rect 32263 10764 32312 10792
rect 32263 10761 32275 10764
rect 32217 10755 32275 10761
rect 32306 10752 32312 10764
rect 32364 10752 32370 10804
rect 32582 10752 32588 10804
rect 32640 10752 32646 10804
rect 33686 10752 33692 10804
rect 33744 10752 33750 10804
rect 35069 10795 35127 10801
rect 35069 10761 35081 10795
rect 35115 10792 35127 10795
rect 35618 10792 35624 10804
rect 35115 10764 35624 10792
rect 35115 10761 35127 10764
rect 35069 10755 35127 10761
rect 35618 10752 35624 10764
rect 35676 10752 35682 10804
rect 28537 10727 28595 10733
rect 28537 10693 28549 10727
rect 28583 10724 28595 10727
rect 28583 10696 28856 10724
rect 28583 10693 28595 10696
rect 28537 10687 28595 10693
rect 28828 10668 28856 10696
rect 29086 10684 29092 10736
rect 29144 10724 29150 10736
rect 32600 10724 32628 10752
rect 29144 10696 30512 10724
rect 29144 10684 29150 10696
rect 28261 10659 28319 10665
rect 28261 10625 28273 10659
rect 28307 10625 28319 10659
rect 28261 10619 28319 10625
rect 28350 10616 28356 10668
rect 28408 10656 28414 10668
rect 28721 10659 28779 10665
rect 28721 10656 28733 10659
rect 28408 10628 28733 10656
rect 28408 10616 28414 10628
rect 28721 10625 28733 10628
rect 28767 10625 28779 10659
rect 28721 10619 28779 10625
rect 28810 10616 28816 10668
rect 28868 10616 28874 10668
rect 28905 10659 28963 10665
rect 28905 10625 28917 10659
rect 28951 10656 28963 10659
rect 28994 10656 29000 10668
rect 28951 10628 29000 10656
rect 28951 10625 28963 10628
rect 28905 10619 28963 10625
rect 28994 10616 29000 10628
rect 29052 10616 29058 10668
rect 30282 10616 30288 10668
rect 30340 10616 30346 10668
rect 30484 10665 30512 10696
rect 32324 10696 32628 10724
rect 30469 10659 30527 10665
rect 30469 10625 30481 10659
rect 30515 10656 30527 10659
rect 31846 10656 31852 10668
rect 30515 10628 31852 10656
rect 30515 10625 30527 10628
rect 30469 10619 30527 10625
rect 31846 10616 31852 10628
rect 31904 10616 31910 10668
rect 32125 10659 32183 10665
rect 32125 10625 32137 10659
rect 32171 10656 32183 10659
rect 32214 10656 32220 10668
rect 32171 10628 32220 10656
rect 32171 10625 32183 10628
rect 32125 10619 32183 10625
rect 32214 10616 32220 10628
rect 32272 10616 32278 10668
rect 32324 10665 32352 10696
rect 32309 10659 32367 10665
rect 32309 10625 32321 10659
rect 32355 10625 32367 10659
rect 32309 10619 32367 10625
rect 32585 10659 32643 10665
rect 32585 10625 32597 10659
rect 32631 10656 32643 10659
rect 32766 10656 32772 10668
rect 32631 10628 32772 10656
rect 32631 10625 32643 10628
rect 32585 10619 32643 10625
rect 32766 10616 32772 10628
rect 32824 10616 32830 10668
rect 33502 10616 33508 10668
rect 33560 10616 33566 10668
rect 33781 10659 33839 10665
rect 33781 10625 33793 10659
rect 33827 10625 33839 10659
rect 33781 10619 33839 10625
rect 34057 10659 34115 10665
rect 34057 10625 34069 10659
rect 34103 10625 34115 10659
rect 34057 10619 34115 10625
rect 23385 10591 23443 10597
rect 23385 10557 23397 10591
rect 23431 10557 23443 10591
rect 23385 10551 23443 10557
rect 23750 10548 23756 10600
rect 23808 10588 23814 10600
rect 23937 10591 23995 10597
rect 23937 10588 23949 10591
rect 23808 10560 23949 10588
rect 23808 10548 23814 10560
rect 23937 10557 23949 10560
rect 23983 10588 23995 10591
rect 24394 10588 24400 10600
rect 23983 10560 24400 10588
rect 23983 10557 23995 10560
rect 23937 10551 23995 10557
rect 24394 10548 24400 10560
rect 24452 10548 24458 10600
rect 30377 10591 30435 10597
rect 24596 10560 28856 10588
rect 24596 10529 24624 10560
rect 24581 10523 24639 10529
rect 21876 10492 22048 10520
rect 22112 10492 24072 10520
rect 21876 10480 21882 10492
rect 17034 10452 17040 10464
rect 10980 10424 17040 10452
rect 10597 10415 10655 10421
rect 17034 10412 17040 10424
rect 17092 10412 17098 10464
rect 18046 10412 18052 10464
rect 18104 10412 18110 10464
rect 20162 10412 20168 10464
rect 20220 10412 20226 10464
rect 20993 10455 21051 10461
rect 20993 10421 21005 10455
rect 21039 10452 21051 10455
rect 21082 10452 21088 10464
rect 21039 10424 21088 10452
rect 21039 10421 21051 10424
rect 20993 10415 21051 10421
rect 21082 10412 21088 10424
rect 21140 10412 21146 10464
rect 21177 10455 21235 10461
rect 21177 10421 21189 10455
rect 21223 10452 21235 10455
rect 21634 10452 21640 10464
rect 21223 10424 21640 10452
rect 21223 10421 21235 10424
rect 21177 10415 21235 10421
rect 21634 10412 21640 10424
rect 21692 10412 21698 10464
rect 22020 10452 22048 10492
rect 24044 10464 24072 10492
rect 24581 10489 24593 10523
rect 24627 10489 24639 10523
rect 28166 10520 28172 10532
rect 24581 10483 24639 10489
rect 27632 10492 28172 10520
rect 22370 10452 22376 10464
rect 22020 10424 22376 10452
rect 22370 10412 22376 10424
rect 22428 10412 22434 10464
rect 22738 10412 22744 10464
rect 22796 10412 22802 10464
rect 24026 10412 24032 10464
rect 24084 10412 24090 10464
rect 27632 10461 27660 10492
rect 28166 10480 28172 10492
rect 28224 10480 28230 10532
rect 28721 10523 28779 10529
rect 28721 10489 28733 10523
rect 28767 10489 28779 10523
rect 28828 10520 28856 10560
rect 30377 10557 30389 10591
rect 30423 10588 30435 10591
rect 32490 10588 32496 10600
rect 30423 10560 32496 10588
rect 30423 10557 30435 10560
rect 30377 10551 30435 10557
rect 32490 10548 32496 10560
rect 32548 10548 32554 10600
rect 32599 10560 32904 10588
rect 32599 10520 32627 10560
rect 28828 10492 32627 10520
rect 32876 10520 32904 10560
rect 33226 10548 33232 10600
rect 33284 10588 33290 10600
rect 33796 10588 33824 10619
rect 33284 10560 33824 10588
rect 33965 10591 34023 10597
rect 33284 10548 33290 10560
rect 33965 10557 33977 10591
rect 34011 10557 34023 10591
rect 33965 10551 34023 10557
rect 33980 10520 34008 10551
rect 32876 10492 34008 10520
rect 28721 10483 28779 10489
rect 27617 10455 27675 10461
rect 27617 10421 27629 10455
rect 27663 10421 27675 10455
rect 27617 10415 27675 10421
rect 27890 10412 27896 10464
rect 27948 10452 27954 10464
rect 28736 10452 28764 10483
rect 32122 10452 32128 10464
rect 27948 10424 32128 10452
rect 27948 10412 27954 10424
rect 32122 10412 32128 10424
rect 32180 10412 32186 10464
rect 32858 10412 32864 10464
rect 32916 10412 32922 10464
rect 33505 10455 33563 10461
rect 33505 10421 33517 10455
rect 33551 10452 33563 10455
rect 34072 10452 34100 10619
rect 34422 10616 34428 10668
rect 34480 10656 34486 10668
rect 34701 10659 34759 10665
rect 34701 10656 34713 10659
rect 34480 10628 34713 10656
rect 34480 10616 34486 10628
rect 34701 10625 34713 10628
rect 34747 10625 34759 10659
rect 34701 10619 34759 10625
rect 34609 10591 34667 10597
rect 34609 10557 34621 10591
rect 34655 10557 34667 10591
rect 34609 10551 34667 10557
rect 34425 10523 34483 10529
rect 34425 10489 34437 10523
rect 34471 10520 34483 10523
rect 34624 10520 34652 10551
rect 34471 10492 34652 10520
rect 34471 10489 34483 10492
rect 34425 10483 34483 10489
rect 33551 10424 34100 10452
rect 33551 10421 33563 10424
rect 33505 10415 33563 10421
rect 1104 10362 38272 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38272 10362
rect 1104 10288 38272 10310
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 4706 10248 4712 10260
rect 4663 10220 4712 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 6178 10208 6184 10260
rect 6236 10208 6242 10260
rect 6362 10208 6368 10260
rect 6420 10208 6426 10260
rect 7558 10208 7564 10260
rect 7616 10248 7622 10260
rect 9950 10248 9956 10260
rect 7616 10220 9956 10248
rect 7616 10208 7622 10220
rect 9950 10208 9956 10220
rect 10008 10248 10014 10260
rect 10008 10220 10732 10248
rect 10008 10208 10014 10220
rect 6380 10180 6408 10208
rect 10704 10192 10732 10220
rect 11790 10208 11796 10260
rect 11848 10248 11854 10260
rect 12158 10248 12164 10260
rect 11848 10220 12164 10248
rect 11848 10208 11854 10220
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 13078 10248 13084 10260
rect 12400 10220 13084 10248
rect 12400 10208 12406 10220
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 14366 10248 14372 10260
rect 13964 10220 14372 10248
rect 13964 10208 13970 10220
rect 14366 10208 14372 10220
rect 14424 10248 14430 10260
rect 17126 10248 17132 10260
rect 14424 10220 17132 10248
rect 14424 10208 14430 10220
rect 17126 10208 17132 10220
rect 17184 10208 17190 10260
rect 18690 10248 18696 10260
rect 17604 10220 18696 10248
rect 8018 10180 8024 10192
rect 5644 10152 6408 10180
rect 7668 10152 8024 10180
rect 5644 10121 5672 10152
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 5810 10072 5816 10124
rect 5868 10072 5874 10124
rect 5902 10072 5908 10124
rect 5960 10112 5966 10124
rect 5960 10084 6224 10112
rect 5960 10072 5966 10084
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10044 3019 10047
rect 3142 10044 3148 10056
rect 3007 10016 3148 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3326 10004 3332 10056
rect 3384 10004 3390 10056
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10044 4859 10047
rect 5537 10047 5595 10053
rect 4847 10016 5212 10044
rect 4847 10013 4859 10016
rect 4801 10007 4859 10013
rect 2777 9979 2835 9985
rect 2777 9945 2789 9979
rect 2823 9976 2835 9979
rect 3344 9976 3372 10004
rect 2823 9948 3372 9976
rect 2823 9945 2835 9948
rect 2777 9939 2835 9945
rect 3142 9868 3148 9920
rect 3200 9868 3206 9920
rect 5184 9917 5212 10016
rect 5537 10013 5549 10047
rect 5583 10044 5595 10047
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5583 10016 6009 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 5997 10013 6009 10016
rect 6043 10044 6055 10047
rect 6086 10044 6092 10056
rect 6043 10016 6092 10044
rect 6043 10013 6055 10016
rect 5997 10007 6055 10013
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 6196 10053 6224 10084
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 7466 10004 7472 10056
rect 7524 10004 7530 10056
rect 7668 10044 7696 10152
rect 8018 10140 8024 10152
rect 8076 10140 8082 10192
rect 8481 10183 8539 10189
rect 8481 10149 8493 10183
rect 8527 10180 8539 10183
rect 9490 10180 9496 10192
rect 8527 10152 9076 10180
rect 8527 10149 8539 10152
rect 8481 10143 8539 10149
rect 7745 10115 7803 10121
rect 7745 10081 7757 10115
rect 7791 10112 7803 10115
rect 8202 10112 8208 10124
rect 7791 10084 8208 10112
rect 7791 10081 7803 10084
rect 7745 10075 7803 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 8322 10115 8380 10121
rect 8322 10081 8334 10115
rect 8368 10112 8380 10115
rect 8662 10112 8668 10124
rect 8368 10084 8668 10112
rect 8368 10081 8380 10084
rect 8322 10075 8380 10081
rect 8662 10072 8668 10084
rect 8720 10072 8726 10124
rect 9048 10121 9076 10152
rect 9232 10152 9496 10180
rect 9033 10115 9091 10121
rect 9033 10081 9045 10115
rect 9079 10081 9091 10115
rect 9033 10075 9091 10081
rect 7837 10047 7895 10053
rect 7837 10044 7849 10047
rect 7668 10016 7849 10044
rect 7837 10013 7849 10016
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 7984 10016 8248 10044
rect 7984 10004 7990 10016
rect 8220 9917 8248 10016
rect 8938 10004 8944 10056
rect 8996 10044 9002 10056
rect 9232 10053 9260 10152
rect 9490 10140 9496 10152
rect 9548 10140 9554 10192
rect 10686 10140 10692 10192
rect 10744 10140 10750 10192
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10112 9367 10115
rect 9766 10112 9772 10124
rect 9355 10084 9772 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 11701 10115 11759 10121
rect 11701 10081 11713 10115
rect 11747 10112 11759 10115
rect 11808 10112 11836 10208
rect 17604 10121 17632 10220
rect 18690 10208 18696 10220
rect 18748 10248 18754 10260
rect 19242 10248 19248 10260
rect 18748 10220 19248 10248
rect 18748 10208 18754 10220
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 20254 10208 20260 10260
rect 20312 10208 20318 10260
rect 20441 10251 20499 10257
rect 20441 10217 20453 10251
rect 20487 10248 20499 10251
rect 20901 10251 20959 10257
rect 20487 10220 20760 10248
rect 20487 10217 20499 10220
rect 20441 10211 20499 10217
rect 11747 10084 11836 10112
rect 17589 10115 17647 10121
rect 11747 10081 11759 10084
rect 11701 10075 11759 10081
rect 17589 10081 17601 10115
rect 17635 10081 17647 10115
rect 20272 10112 20300 10208
rect 20530 10140 20536 10192
rect 20588 10180 20594 10192
rect 20588 10152 20684 10180
rect 20588 10140 20594 10152
rect 17589 10075 17647 10081
rect 18340 10084 18828 10112
rect 20272 10084 20576 10112
rect 18340 10056 18368 10084
rect 18800 10056 18828 10084
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 8996 10016 9137 10044
rect 8996 10004 9002 10016
rect 9125 10013 9137 10016
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 8478 9936 8484 9988
rect 8536 9976 8542 9988
rect 9232 9976 9260 10007
rect 11422 10004 11428 10056
rect 11480 10004 11486 10056
rect 13262 10004 13268 10056
rect 13320 10004 13326 10056
rect 13722 10004 13728 10056
rect 13780 10004 13786 10056
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10013 17831 10047
rect 17773 10007 17831 10013
rect 11977 9979 12035 9985
rect 11977 9976 11989 9979
rect 8536 9948 9260 9976
rect 11624 9948 11989 9976
rect 8536 9936 8542 9948
rect 5169 9911 5227 9917
rect 5169 9877 5181 9911
rect 5215 9877 5227 9911
rect 5169 9871 5227 9877
rect 7745 9911 7803 9917
rect 7745 9877 7757 9911
rect 7791 9908 7803 9911
rect 8113 9911 8171 9917
rect 8113 9908 8125 9911
rect 7791 9880 8125 9908
rect 7791 9877 7803 9880
rect 7745 9871 7803 9877
rect 8113 9877 8125 9880
rect 8159 9877 8171 9911
rect 8113 9871 8171 9877
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 9490 9868 9496 9920
rect 9548 9868 9554 9920
rect 11624 9917 11652 9948
rect 11977 9945 11989 9948
rect 12023 9945 12035 9979
rect 13280 9976 13308 10004
rect 17788 9976 17816 10007
rect 18046 10004 18052 10056
rect 18104 10004 18110 10056
rect 18230 10004 18236 10056
rect 18288 10004 18294 10056
rect 18322 10004 18328 10056
rect 18380 10004 18386 10056
rect 18414 10004 18420 10056
rect 18472 10004 18478 10056
rect 18782 10004 18788 10056
rect 18840 10004 18846 10056
rect 20162 10004 20168 10056
rect 20220 10044 20226 10056
rect 20257 10047 20315 10053
rect 20257 10044 20269 10047
rect 20220 10016 20269 10044
rect 20220 10004 20226 10016
rect 20257 10013 20269 10016
rect 20303 10013 20315 10047
rect 20257 10007 20315 10013
rect 20438 10004 20444 10056
rect 20496 10004 20502 10056
rect 20548 10053 20576 10084
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10013 20591 10047
rect 20656 10044 20684 10152
rect 20732 10112 20760 10220
rect 20901 10217 20913 10251
rect 20947 10248 20959 10251
rect 21818 10248 21824 10260
rect 20947 10220 21824 10248
rect 20947 10217 20959 10220
rect 20901 10211 20959 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 22370 10208 22376 10260
rect 22428 10208 22434 10260
rect 22462 10208 22468 10260
rect 22520 10248 22526 10260
rect 22649 10251 22707 10257
rect 22649 10248 22661 10251
rect 22520 10220 22661 10248
rect 22520 10208 22526 10220
rect 22649 10217 22661 10220
rect 22695 10217 22707 10251
rect 22649 10211 22707 10217
rect 22738 10208 22744 10260
rect 22796 10208 22802 10260
rect 25682 10208 25688 10260
rect 25740 10248 25746 10260
rect 28442 10248 28448 10260
rect 25740 10220 28448 10248
rect 25740 10208 25746 10220
rect 28442 10208 28448 10220
rect 28500 10248 28506 10260
rect 28500 10220 29316 10248
rect 28500 10208 28506 10220
rect 20809 10183 20867 10189
rect 20809 10149 20821 10183
rect 20855 10180 20867 10183
rect 21177 10183 21235 10189
rect 21177 10180 21189 10183
rect 20855 10152 21189 10180
rect 20855 10149 20867 10152
rect 20809 10143 20867 10149
rect 21177 10149 21189 10152
rect 21223 10149 21235 10183
rect 21637 10183 21695 10189
rect 21637 10180 21649 10183
rect 21177 10143 21235 10149
rect 21376 10152 21649 10180
rect 21376 10121 21404 10152
rect 21637 10149 21649 10152
rect 21683 10149 21695 10183
rect 21637 10143 21695 10149
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 20732 10084 21281 10112
rect 21269 10081 21281 10084
rect 21315 10081 21327 10115
rect 21269 10075 21327 10081
rect 21361 10115 21419 10121
rect 21361 10081 21373 10115
rect 21407 10081 21419 10115
rect 22373 10115 22431 10121
rect 21361 10075 21419 10081
rect 21560 10084 22232 10112
rect 21085 10047 21143 10053
rect 20656 10016 21052 10044
rect 20533 10007 20591 10013
rect 11977 9939 12035 9945
rect 12406 9948 12466 9976
rect 13280 9948 17816 9976
rect 17957 9979 18015 9985
rect 11609 9911 11667 9917
rect 11609 9877 11621 9911
rect 11655 9877 11667 9911
rect 11609 9871 11667 9877
rect 12158 9868 12164 9920
rect 12216 9908 12222 9920
rect 12406 9908 12434 9948
rect 17957 9945 17969 9979
rect 18003 9976 18015 9979
rect 19337 9979 19395 9985
rect 19337 9976 19349 9979
rect 18003 9948 19349 9976
rect 18003 9945 18015 9948
rect 17957 9939 18015 9945
rect 19337 9945 19349 9948
rect 19383 9945 19395 9979
rect 19337 9939 19395 9945
rect 19705 9979 19763 9985
rect 19705 9945 19717 9979
rect 19751 9976 19763 9979
rect 20346 9976 20352 9988
rect 19751 9948 20352 9976
rect 19751 9945 19763 9948
rect 19705 9939 19763 9945
rect 20346 9936 20352 9948
rect 20404 9936 20410 9988
rect 20622 9936 20628 9988
rect 20680 9936 20686 9988
rect 20809 9979 20867 9985
rect 20809 9945 20821 9979
rect 20855 9976 20867 9979
rect 20898 9976 20904 9988
rect 20855 9948 20904 9976
rect 20855 9945 20867 9948
rect 20809 9939 20867 9945
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 21024 9976 21052 10016
rect 21085 10013 21097 10047
rect 21131 10044 21143 10047
rect 21174 10044 21180 10056
rect 21131 10016 21180 10044
rect 21131 10013 21143 10016
rect 21085 10007 21143 10013
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 21560 10053 21588 10084
rect 22204 10056 22232 10084
rect 22373 10081 22385 10115
rect 22419 10112 22431 10115
rect 22756 10112 22784 10208
rect 24118 10140 24124 10192
rect 24176 10180 24182 10192
rect 28902 10180 28908 10192
rect 24176 10152 28908 10180
rect 24176 10140 24182 10152
rect 28902 10140 28908 10152
rect 28960 10140 28966 10192
rect 28997 10183 29055 10189
rect 28997 10149 29009 10183
rect 29043 10180 29055 10183
rect 29086 10180 29092 10192
rect 29043 10152 29092 10180
rect 29043 10149 29055 10152
rect 28997 10143 29055 10149
rect 29086 10140 29092 10152
rect 29144 10140 29150 10192
rect 29288 10180 29316 10220
rect 30742 10208 30748 10260
rect 30800 10208 30806 10260
rect 32677 10251 32735 10257
rect 32677 10217 32689 10251
rect 32723 10248 32735 10251
rect 32766 10248 32772 10260
rect 32723 10220 32772 10248
rect 32723 10217 32735 10220
rect 32677 10211 32735 10217
rect 32766 10208 32772 10220
rect 32824 10208 32830 10260
rect 33502 10208 33508 10260
rect 33560 10208 33566 10260
rect 30760 10180 30788 10208
rect 32950 10180 32956 10192
rect 29288 10152 30788 10180
rect 32600 10152 32956 10180
rect 22419 10084 22784 10112
rect 22419 10081 22431 10084
rect 22373 10075 22431 10081
rect 26418 10072 26424 10124
rect 26476 10112 26482 10124
rect 27890 10112 27896 10124
rect 26476 10084 27896 10112
rect 26476 10072 26482 10084
rect 27890 10072 27896 10084
rect 27948 10072 27954 10124
rect 28166 10072 28172 10124
rect 28224 10112 28230 10124
rect 28224 10084 30144 10112
rect 28224 10072 28230 10084
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10013 21603 10047
rect 21545 10007 21603 10013
rect 21634 10004 21640 10056
rect 21692 10004 21698 10056
rect 21818 10004 21824 10056
rect 21876 10004 21882 10056
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10013 21971 10047
rect 21913 10007 21971 10013
rect 21928 9976 21956 10007
rect 22186 10004 22192 10056
rect 22244 10004 22250 10056
rect 22278 10004 22284 10056
rect 22336 10004 22342 10056
rect 22554 10004 22560 10056
rect 22612 10044 22618 10056
rect 26142 10044 26148 10056
rect 22612 10016 26148 10044
rect 22612 10004 22618 10016
rect 26142 10004 26148 10016
rect 26200 10004 26206 10056
rect 28261 10047 28319 10053
rect 28261 10044 28273 10047
rect 27908 10016 28273 10044
rect 27908 9988 27936 10016
rect 28261 10013 28273 10016
rect 28307 10013 28319 10047
rect 28261 10007 28319 10013
rect 28350 10004 28356 10056
rect 28408 10044 28414 10056
rect 28629 10047 28687 10053
rect 28629 10044 28641 10047
rect 28408 10016 28641 10044
rect 28408 10004 28414 10016
rect 28629 10013 28641 10016
rect 28675 10013 28687 10047
rect 28629 10007 28687 10013
rect 28718 10004 28724 10056
rect 28776 10004 28782 10056
rect 28902 10004 28908 10056
rect 28960 10004 28966 10056
rect 30116 10053 30144 10084
rect 30374 10072 30380 10124
rect 30432 10072 30438 10124
rect 30484 10121 30512 10152
rect 30469 10115 30527 10121
rect 30469 10081 30481 10115
rect 30515 10081 30527 10115
rect 30469 10075 30527 10081
rect 30101 10047 30159 10053
rect 30101 10013 30113 10047
rect 30147 10013 30159 10047
rect 30101 10007 30159 10013
rect 30190 10004 30196 10056
rect 30248 10042 30254 10056
rect 30285 10047 30343 10053
rect 30285 10042 30297 10047
rect 30248 10014 30297 10042
rect 30248 10004 30254 10014
rect 30285 10013 30297 10014
rect 30331 10013 30343 10047
rect 30285 10007 30343 10013
rect 30650 10004 30656 10056
rect 30708 10044 30714 10056
rect 32600 10053 32628 10152
rect 32950 10140 32956 10152
rect 33008 10140 33014 10192
rect 32876 10084 33916 10112
rect 32876 10056 32904 10084
rect 32585 10047 32643 10053
rect 32585 10044 32597 10047
rect 30708 10016 32597 10044
rect 30708 10004 30714 10016
rect 32585 10013 32597 10016
rect 32631 10013 32643 10047
rect 32585 10007 32643 10013
rect 32858 10004 32864 10056
rect 32916 10004 32922 10056
rect 33888 10053 33916 10084
rect 33781 10047 33839 10053
rect 33781 10013 33793 10047
rect 33827 10013 33839 10047
rect 33781 10007 33839 10013
rect 33873 10047 33931 10053
rect 33873 10013 33885 10047
rect 33919 10013 33931 10047
rect 33873 10007 33931 10013
rect 26326 9976 26332 9988
rect 21024 9948 21956 9976
rect 22204 9948 26332 9976
rect 12216 9880 12434 9908
rect 12216 9868 12222 9880
rect 13446 9868 13452 9920
rect 13504 9908 13510 9920
rect 16666 9908 16672 9920
rect 13504 9880 16672 9908
rect 13504 9868 13510 9880
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 18693 9911 18751 9917
rect 18693 9877 18705 9911
rect 18739 9908 18751 9911
rect 22204 9908 22232 9948
rect 26326 9936 26332 9948
rect 26384 9936 26390 9988
rect 27890 9936 27896 9988
rect 27948 9936 27954 9988
rect 28445 9979 28503 9985
rect 28445 9945 28457 9979
rect 28491 9976 28503 9979
rect 28994 9976 29000 9988
rect 28491 9948 29000 9976
rect 28491 9945 28503 9948
rect 28445 9939 28503 9945
rect 28994 9936 29000 9948
rect 29052 9976 29058 9988
rect 33796 9976 33824 10007
rect 33962 10004 33968 10056
rect 34020 10004 34026 10056
rect 34054 10004 34060 10056
rect 34112 10044 34118 10056
rect 34149 10047 34207 10053
rect 34149 10044 34161 10047
rect 34112 10016 34161 10044
rect 34112 10004 34118 10016
rect 34149 10013 34161 10016
rect 34195 10013 34207 10047
rect 34149 10007 34207 10013
rect 29052 9948 33824 9976
rect 29052 9936 29058 9948
rect 18739 9880 22232 9908
rect 18739 9877 18751 9880
rect 18693 9871 18751 9877
rect 22922 9868 22928 9920
rect 22980 9908 22986 9920
rect 24854 9908 24860 9920
rect 22980 9880 24860 9908
rect 22980 9868 22986 9880
rect 24854 9868 24860 9880
rect 24912 9868 24918 9920
rect 24946 9868 24952 9920
rect 25004 9908 25010 9920
rect 28902 9908 28908 9920
rect 25004 9880 28908 9908
rect 25004 9868 25010 9880
rect 28902 9868 28908 9880
rect 28960 9868 28966 9920
rect 30834 9868 30840 9920
rect 30892 9868 30898 9920
rect 1104 9818 38272 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38272 9818
rect 1104 9744 38272 9766
rect 3142 9664 3148 9716
rect 3200 9664 3206 9716
rect 8128 9676 8708 9704
rect 3160 9636 3188 9664
rect 3160 9608 3464 9636
rect 3234 9528 3240 9580
rect 3292 9528 3298 9580
rect 3436 9577 3464 9608
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 6365 9639 6423 9645
rect 6365 9636 6377 9639
rect 5592 9608 6377 9636
rect 5592 9596 5598 9608
rect 6365 9605 6377 9608
rect 6411 9605 6423 9639
rect 8128 9636 8156 9676
rect 6365 9599 6423 9605
rect 6748 9608 8156 9636
rect 6748 9580 6776 9608
rect 8202 9596 8208 9648
rect 8260 9636 8266 9648
rect 8297 9639 8355 9645
rect 8297 9636 8309 9639
rect 8260 9608 8309 9636
rect 8260 9596 8266 9608
rect 8297 9605 8309 9608
rect 8343 9636 8355 9639
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 8343 9608 8585 9636
rect 8343 9605 8355 9608
rect 8297 9599 8355 9605
rect 8573 9605 8585 9608
rect 8619 9605 8631 9639
rect 8680 9636 8708 9676
rect 11422 9664 11428 9716
rect 11480 9704 11486 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11480 9676 11805 9704
rect 11480 9664 11486 9676
rect 11793 9673 11805 9676
rect 11839 9673 11851 9707
rect 11793 9667 11851 9673
rect 13078 9664 13084 9716
rect 13136 9664 13142 9716
rect 13446 9664 13452 9716
rect 13504 9664 13510 9716
rect 15933 9707 15991 9713
rect 15212 9676 15608 9704
rect 10594 9636 10600 9648
rect 8680 9608 10600 9636
rect 8573 9599 8631 9605
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 10781 9639 10839 9645
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 11606 9636 11612 9648
rect 10827 9608 11612 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 11606 9596 11612 9608
rect 11664 9596 11670 9648
rect 11698 9596 11704 9648
rect 11756 9636 11762 9648
rect 13170 9636 13176 9648
rect 11756 9608 13176 9636
rect 11756 9596 11762 9608
rect 13170 9596 13176 9608
rect 13228 9596 13234 9648
rect 14366 9636 14372 9648
rect 13280 9608 13768 9636
rect 3329 9571 3387 9577
rect 3329 9537 3341 9571
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9568 3663 9571
rect 3694 9568 3700 9580
rect 3651 9540 3700 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 3344 9500 3372 9531
rect 3694 9528 3700 9540
rect 3752 9568 3758 9580
rect 6641 9571 6699 9577
rect 3752 9540 4752 9568
rect 3752 9528 3758 9540
rect 3344 9472 4016 9500
rect 3988 9376 4016 9472
rect 4724 9376 4752 9540
rect 6641 9537 6653 9571
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 6656 9500 6684 9531
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 6822 9528 6828 9580
rect 6880 9528 6886 9580
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9568 7067 9571
rect 7098 9568 7104 9580
rect 7055 9540 7104 9568
rect 7055 9537 7067 9540
rect 7009 9531 7067 9537
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 7834 9568 7840 9580
rect 7791 9540 7840 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8110 9568 8116 9580
rect 8067 9540 8116 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8110 9528 8116 9540
rect 8168 9528 8174 9580
rect 8478 9528 8484 9580
rect 8536 9528 8542 9580
rect 8665 9571 8723 9577
rect 8665 9537 8677 9571
rect 8711 9568 8723 9571
rect 8938 9568 8944 9580
rect 8711 9540 8944 9568
rect 8711 9537 8723 9540
rect 8665 9531 8723 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9568 10287 9571
rect 10275 9540 10364 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 6656 9472 9536 9500
rect 7466 9392 7472 9444
rect 7524 9392 7530 9444
rect 8021 9435 8079 9441
rect 8021 9401 8033 9435
rect 8067 9432 8079 9435
rect 8202 9432 8208 9444
rect 8067 9404 8208 9432
rect 8067 9401 8079 9404
rect 8021 9395 8079 9401
rect 8202 9392 8208 9404
rect 8260 9392 8266 9444
rect 9508 9432 9536 9472
rect 10336 9441 10364 9540
rect 10686 9528 10692 9580
rect 10744 9568 10750 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 10744 9540 12173 9568
rect 10744 9528 10750 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9568 12311 9571
rect 13280 9568 13308 9608
rect 13740 9580 13768 9608
rect 13832 9608 14372 9636
rect 13832 9580 13860 9608
rect 14366 9596 14372 9608
rect 14424 9596 14430 9648
rect 12299 9540 13308 9568
rect 12299 9537 12311 9540
rect 12253 9531 12311 9537
rect 13722 9528 13728 9580
rect 13780 9528 13786 9580
rect 13814 9528 13820 9580
rect 13872 9528 13878 9580
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 15212 9568 15240 9676
rect 15286 9596 15292 9648
rect 15344 9636 15350 9648
rect 15473 9639 15531 9645
rect 15473 9636 15485 9639
rect 15344 9608 15485 9636
rect 15344 9596 15350 9608
rect 15473 9605 15485 9608
rect 15519 9605 15531 9639
rect 15580 9636 15608 9676
rect 15933 9673 15945 9707
rect 15979 9673 15991 9707
rect 15933 9667 15991 9673
rect 15580 9608 15884 9636
rect 15473 9599 15531 9605
rect 14148 9540 15240 9568
rect 14148 9528 14154 9540
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 15565 9571 15623 9577
rect 15565 9568 15577 9571
rect 15436 9540 15577 9568
rect 15436 9528 15442 9540
rect 15565 9537 15577 9540
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 10870 9460 10876 9512
rect 10928 9460 10934 9512
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9500 12495 9503
rect 12618 9500 12624 9512
rect 12483 9472 12624 9500
rect 12483 9469 12495 9472
rect 12437 9463 12495 9469
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 13262 9460 13268 9512
rect 13320 9500 13326 9512
rect 13541 9503 13599 9509
rect 13541 9500 13553 9503
rect 13320 9472 13553 9500
rect 13320 9460 13326 9472
rect 13541 9469 13553 9472
rect 13587 9469 13599 9503
rect 13541 9463 13599 9469
rect 13633 9503 13691 9509
rect 13633 9469 13645 9503
rect 13679 9500 13691 9503
rect 15194 9500 15200 9512
rect 13679 9472 15200 9500
rect 13679 9469 13691 9472
rect 13633 9463 13691 9469
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 15289 9503 15347 9509
rect 15289 9469 15301 9503
rect 15335 9500 15347 9503
rect 15654 9500 15660 9512
rect 15335 9472 15660 9500
rect 15335 9469 15347 9472
rect 15289 9463 15347 9469
rect 15654 9460 15660 9472
rect 15712 9460 15718 9512
rect 15856 9500 15884 9608
rect 15948 9568 15976 9667
rect 20254 9664 20260 9716
rect 20312 9664 20318 9716
rect 22370 9664 22376 9716
rect 22428 9704 22434 9716
rect 22465 9707 22523 9713
rect 22465 9704 22477 9707
rect 22428 9676 22477 9704
rect 22428 9664 22434 9676
rect 22465 9673 22477 9676
rect 22511 9673 22523 9707
rect 23014 9704 23020 9716
rect 22465 9667 22523 9673
rect 22664 9676 23020 9704
rect 18046 9596 18052 9648
rect 18104 9636 18110 9648
rect 20272 9636 20300 9664
rect 18104 9608 18828 9636
rect 18104 9596 18110 9608
rect 16209 9571 16267 9577
rect 16209 9568 16221 9571
rect 15948 9540 16221 9568
rect 16209 9537 16221 9540
rect 16255 9537 16267 9571
rect 16209 9531 16267 9537
rect 16666 9528 16672 9580
rect 16724 9568 16730 9580
rect 16761 9571 16819 9577
rect 16761 9568 16773 9571
rect 16724 9540 16773 9568
rect 16724 9528 16730 9540
rect 16761 9537 16773 9540
rect 16807 9568 16819 9571
rect 17310 9568 17316 9580
rect 16807 9540 17316 9568
rect 16807 9537 16819 9540
rect 16761 9531 16819 9537
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 18322 9528 18328 9580
rect 18380 9568 18386 9580
rect 18800 9577 18828 9608
rect 19812 9608 20300 9636
rect 19812 9577 19840 9608
rect 18417 9571 18475 9577
rect 18417 9568 18429 9571
rect 18380 9540 18429 9568
rect 18380 9528 18386 9540
rect 18417 9537 18429 9540
rect 18463 9537 18475 9571
rect 18417 9531 18475 9537
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9537 18843 9571
rect 18785 9531 18843 9537
rect 19797 9571 19855 9577
rect 19797 9537 19809 9571
rect 19843 9537 19855 9571
rect 19797 9531 19855 9537
rect 19886 9528 19892 9580
rect 19944 9528 19950 9580
rect 20073 9571 20131 9577
rect 20073 9537 20085 9571
rect 20119 9568 20131 9571
rect 20162 9568 20168 9580
rect 20119 9540 20168 9568
rect 20119 9537 20131 9540
rect 20073 9531 20131 9537
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 22664 9577 22692 9676
rect 23014 9664 23020 9676
rect 23072 9704 23078 9716
rect 23474 9704 23480 9716
rect 23072 9676 23480 9704
rect 23072 9664 23078 9676
rect 23474 9664 23480 9676
rect 23532 9664 23538 9716
rect 23566 9664 23572 9716
rect 23624 9704 23630 9716
rect 23624 9676 24072 9704
rect 23624 9664 23630 9676
rect 23109 9639 23167 9645
rect 23109 9605 23121 9639
rect 23155 9636 23167 9639
rect 23750 9636 23756 9648
rect 23155 9608 23756 9636
rect 23155 9605 23167 9608
rect 23109 9599 23167 9605
rect 23750 9596 23756 9608
rect 23808 9596 23814 9648
rect 24044 9636 24072 9676
rect 24118 9664 24124 9716
rect 24176 9704 24182 9716
rect 24854 9704 24860 9716
rect 24176 9676 24532 9704
rect 24176 9664 24182 9676
rect 24504 9636 24532 9676
rect 24596 9676 24860 9704
rect 24596 9645 24624 9676
rect 24854 9664 24860 9676
rect 24912 9664 24918 9716
rect 27338 9664 27344 9716
rect 27396 9704 27402 9716
rect 27396 9676 27844 9704
rect 27396 9664 27402 9676
rect 24044 9608 24348 9636
rect 22649 9571 22707 9577
rect 22649 9568 22661 9571
rect 22066 9540 22661 9568
rect 16942 9500 16948 9512
rect 15856 9472 16948 9500
rect 16942 9460 16948 9472
rect 17000 9500 17006 9512
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 17000 9472 17233 9500
rect 17000 9460 17006 9472
rect 17221 9469 17233 9472
rect 17267 9500 17279 9503
rect 17494 9500 17500 9512
rect 17267 9472 17500 9500
rect 17267 9469 17279 9472
rect 17221 9463 17279 9469
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 18230 9460 18236 9512
rect 18288 9460 18294 9512
rect 18693 9503 18751 9509
rect 18693 9500 18705 9503
rect 18432 9472 18705 9500
rect 10321 9435 10379 9441
rect 9508 9404 10272 9432
rect 2958 9324 2964 9376
rect 3016 9324 3022 9376
rect 3970 9324 3976 9376
rect 4028 9324 4034 9376
rect 4706 9324 4712 9376
rect 4764 9324 4770 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 9674 9364 9680 9376
rect 7340 9336 9680 9364
rect 7340 9324 7346 9336
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10042 9324 10048 9376
rect 10100 9324 10106 9376
rect 10244 9364 10272 9404
rect 10321 9401 10333 9435
rect 10367 9401 10379 9435
rect 10321 9395 10379 9401
rect 11422 9392 11428 9444
rect 11480 9432 11486 9444
rect 12158 9432 12164 9444
rect 11480 9404 12164 9432
rect 11480 9392 11486 9404
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 18322 9432 18328 9444
rect 12268 9404 18328 9432
rect 12268 9364 12296 9404
rect 18322 9392 18328 9404
rect 18380 9392 18386 9444
rect 10244 9336 12296 9364
rect 13170 9324 13176 9376
rect 13228 9364 13234 9376
rect 13906 9364 13912 9376
rect 13228 9336 13912 9364
rect 13228 9324 13234 9336
rect 13906 9324 13912 9336
rect 13964 9324 13970 9376
rect 16022 9324 16028 9376
rect 16080 9324 16086 9376
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 18432 9364 18460 9472
rect 18693 9469 18705 9472
rect 18739 9469 18751 9503
rect 18693 9463 18751 9469
rect 19426 9460 19432 9512
rect 19484 9460 19490 9512
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9500 20039 9503
rect 20254 9500 20260 9512
rect 20027 9472 20260 9500
rect 20027 9469 20039 9472
rect 19981 9463 20039 9469
rect 20254 9460 20260 9472
rect 20312 9500 20318 9512
rect 22066 9500 22094 9540
rect 22649 9537 22661 9540
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 22741 9571 22799 9577
rect 22741 9537 22753 9571
rect 22787 9568 22799 9571
rect 23017 9571 23075 9577
rect 22787 9540 22968 9568
rect 22787 9537 22799 9540
rect 22741 9531 22799 9537
rect 20312 9472 22094 9500
rect 20312 9460 20318 9472
rect 19058 9392 19064 9444
rect 19116 9432 19122 9444
rect 22278 9432 22284 9444
rect 19116 9404 22284 9432
rect 19116 9392 19122 9404
rect 22278 9392 22284 9404
rect 22336 9432 22342 9444
rect 22738 9432 22744 9444
rect 22336 9404 22744 9432
rect 22336 9392 22342 9404
rect 22738 9392 22744 9404
rect 22796 9392 22802 9444
rect 16356 9336 18460 9364
rect 16356 9324 16362 9336
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 19613 9367 19671 9373
rect 19613 9364 19625 9367
rect 19392 9336 19625 9364
rect 19392 9324 19398 9336
rect 19613 9333 19625 9336
rect 19659 9333 19671 9367
rect 19613 9327 19671 9333
rect 22554 9324 22560 9376
rect 22612 9364 22618 9376
rect 22940 9364 22968 9540
rect 23017 9537 23029 9571
rect 23063 9568 23075 9571
rect 23063 9540 23336 9568
rect 23063 9537 23075 9540
rect 23017 9531 23075 9537
rect 23308 9512 23336 9540
rect 23382 9528 23388 9580
rect 23440 9568 23446 9580
rect 24320 9577 24348 9608
rect 24412 9608 24532 9636
rect 24581 9639 24639 9645
rect 24412 9577 24440 9608
rect 24581 9605 24593 9639
rect 24627 9605 24639 9639
rect 24581 9599 24639 9605
rect 24673 9639 24731 9645
rect 24673 9605 24685 9639
rect 24719 9636 24731 9639
rect 24946 9636 24952 9648
rect 24719 9608 24952 9636
rect 24719 9605 24731 9608
rect 24673 9599 24731 9605
rect 24946 9596 24952 9608
rect 25004 9596 25010 9648
rect 26329 9639 26387 9645
rect 26329 9605 26341 9639
rect 26375 9636 26387 9639
rect 27816 9636 27844 9676
rect 33134 9664 33140 9716
rect 33192 9704 33198 9716
rect 33229 9707 33287 9713
rect 33229 9704 33241 9707
rect 33192 9676 33241 9704
rect 33192 9664 33198 9676
rect 33229 9673 33241 9676
rect 33275 9704 33287 9707
rect 33962 9704 33968 9716
rect 33275 9676 33968 9704
rect 33275 9673 33287 9676
rect 33229 9667 33287 9673
rect 33962 9664 33968 9676
rect 34020 9664 34026 9716
rect 30009 9639 30067 9645
rect 26375 9608 27752 9636
rect 27816 9608 29960 9636
rect 26375 9605 26387 9608
rect 26329 9599 26387 9605
rect 27724 9580 27752 9608
rect 24121 9574 24179 9577
rect 23952 9571 24179 9574
rect 23952 9568 24133 9571
rect 23440 9546 24133 9568
rect 23440 9540 23980 9546
rect 23440 9528 23446 9540
rect 24121 9537 24133 9546
rect 24167 9537 24179 9571
rect 24121 9531 24179 9537
rect 24305 9571 24363 9577
rect 24305 9537 24317 9571
rect 24351 9537 24363 9571
rect 24305 9531 24363 9537
rect 24397 9571 24455 9577
rect 24397 9537 24409 9571
rect 24443 9537 24455 9571
rect 24765 9571 24823 9577
rect 24765 9568 24777 9571
rect 24397 9531 24455 9537
rect 24688 9540 24777 9568
rect 23290 9460 23296 9512
rect 23348 9460 23354 9512
rect 24320 9500 24348 9531
rect 24688 9500 24716 9540
rect 24765 9537 24777 9540
rect 24811 9537 24823 9571
rect 24765 9531 24823 9537
rect 25961 9571 26019 9577
rect 25961 9537 25973 9571
rect 26007 9537 26019 9571
rect 25961 9531 26019 9537
rect 24320 9472 24716 9500
rect 25498 9460 25504 9512
rect 25556 9500 25562 9512
rect 25976 9500 26004 9531
rect 26142 9528 26148 9580
rect 26200 9568 26206 9580
rect 26421 9571 26479 9577
rect 26421 9568 26433 9571
rect 26200 9540 26433 9568
rect 26200 9528 26206 9540
rect 26421 9537 26433 9540
rect 26467 9537 26479 9571
rect 26421 9531 26479 9537
rect 26605 9571 26663 9577
rect 26605 9537 26617 9571
rect 26651 9537 26663 9571
rect 26605 9531 26663 9537
rect 26973 9571 27031 9577
rect 26973 9537 26985 9571
rect 27019 9537 27031 9571
rect 26973 9531 27031 9537
rect 26620 9500 26648 9531
rect 25556 9472 26648 9500
rect 26988 9500 27016 9531
rect 27062 9528 27068 9580
rect 27120 9568 27126 9580
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 27120 9540 27169 9568
rect 27120 9528 27126 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 27338 9528 27344 9580
rect 27396 9528 27402 9580
rect 27433 9571 27491 9577
rect 27433 9537 27445 9571
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 27356 9500 27384 9528
rect 26988 9472 27384 9500
rect 25556 9460 25562 9472
rect 24302 9392 24308 9444
rect 24360 9392 24366 9444
rect 24949 9435 25007 9441
rect 24949 9401 24961 9435
rect 24995 9432 25007 9435
rect 27448 9432 27476 9531
rect 27706 9528 27712 9580
rect 27764 9528 27770 9580
rect 28718 9528 28724 9580
rect 28776 9568 28782 9580
rect 28813 9571 28871 9577
rect 28813 9568 28825 9571
rect 28776 9540 28825 9568
rect 28776 9528 28782 9540
rect 28813 9537 28825 9540
rect 28859 9537 28871 9571
rect 28813 9531 28871 9537
rect 28902 9528 28908 9580
rect 28960 9568 28966 9580
rect 28997 9571 29055 9577
rect 28997 9568 29009 9571
rect 28960 9540 29009 9568
rect 28960 9528 28966 9540
rect 28997 9537 29009 9540
rect 29043 9537 29055 9571
rect 28997 9531 29055 9537
rect 29638 9528 29644 9580
rect 29696 9528 29702 9580
rect 29730 9528 29736 9580
rect 29788 9528 29794 9580
rect 29932 9577 29960 9608
rect 30009 9605 30021 9639
rect 30055 9636 30067 9639
rect 30055 9608 31754 9636
rect 30055 9605 30067 9608
rect 30009 9599 30067 9605
rect 29825 9571 29883 9577
rect 29825 9537 29837 9571
rect 29871 9537 29883 9571
rect 29825 9531 29883 9537
rect 29917 9571 29975 9577
rect 29917 9537 29929 9571
rect 29963 9537 29975 9571
rect 29917 9531 29975 9537
rect 28736 9432 28764 9528
rect 29840 9500 29868 9531
rect 30098 9528 30104 9580
rect 30156 9528 30162 9580
rect 30742 9528 30748 9580
rect 30800 9528 30806 9580
rect 30834 9528 30840 9580
rect 30892 9568 30898 9580
rect 31021 9571 31079 9577
rect 31021 9568 31033 9571
rect 30892 9540 31033 9568
rect 30892 9528 30898 9540
rect 31021 9537 31033 9540
rect 31067 9537 31079 9571
rect 31021 9531 31079 9537
rect 31297 9571 31355 9577
rect 31297 9537 31309 9571
rect 31343 9568 31355 9571
rect 31386 9568 31392 9580
rect 31343 9540 31392 9568
rect 31343 9537 31355 9540
rect 31297 9531 31355 9537
rect 31386 9528 31392 9540
rect 31444 9528 31450 9580
rect 31573 9571 31631 9577
rect 31573 9537 31585 9571
rect 31619 9537 31631 9571
rect 31573 9531 31631 9537
rect 30190 9500 30196 9512
rect 29840 9472 30196 9500
rect 30190 9460 30196 9472
rect 30248 9460 30254 9512
rect 24995 9404 27476 9432
rect 27540 9404 28764 9432
rect 24995 9401 25007 9404
rect 24949 9395 25007 9401
rect 24118 9364 24124 9376
rect 22612 9336 24124 9364
rect 22612 9324 22618 9336
rect 24118 9324 24124 9336
rect 24176 9324 24182 9376
rect 26510 9324 26516 9376
rect 26568 9364 26574 9376
rect 27540 9364 27568 9404
rect 30926 9392 30932 9444
rect 30984 9432 30990 9444
rect 31205 9435 31263 9441
rect 31205 9432 31217 9435
rect 30984 9404 31217 9432
rect 30984 9392 30990 9404
rect 31205 9401 31217 9404
rect 31251 9401 31263 9435
rect 31205 9395 31263 9401
rect 31588 9376 31616 9531
rect 31726 9500 31754 9608
rect 33042 9596 33048 9648
rect 33100 9596 33106 9648
rect 32493 9571 32551 9577
rect 32493 9537 32505 9571
rect 32539 9568 32551 9571
rect 32766 9568 32772 9580
rect 32539 9540 32772 9568
rect 32539 9537 32551 9540
rect 32493 9531 32551 9537
rect 32766 9528 32772 9540
rect 32824 9528 32830 9580
rect 32861 9571 32919 9577
rect 32861 9537 32873 9571
rect 32907 9537 32919 9571
rect 32861 9531 32919 9537
rect 32401 9503 32459 9509
rect 32401 9500 32413 9503
rect 31726 9472 32413 9500
rect 32401 9469 32413 9472
rect 32447 9469 32459 9503
rect 32401 9463 32459 9469
rect 32030 9392 32036 9444
rect 32088 9432 32094 9444
rect 32125 9435 32183 9441
rect 32125 9432 32137 9435
rect 32088 9404 32137 9432
rect 32088 9392 32094 9404
rect 32125 9401 32137 9404
rect 32171 9432 32183 9435
rect 32876 9432 32904 9531
rect 32171 9404 32904 9432
rect 32171 9401 32183 9404
rect 32125 9395 32183 9401
rect 26568 9336 27568 9364
rect 27617 9367 27675 9373
rect 26568 9324 26574 9336
rect 27617 9333 27629 9367
rect 27663 9364 27675 9367
rect 28074 9364 28080 9376
rect 27663 9336 28080 9364
rect 27663 9333 27675 9336
rect 27617 9327 27675 9333
rect 28074 9324 28080 9336
rect 28132 9324 28138 9376
rect 29181 9367 29239 9373
rect 29181 9333 29193 9367
rect 29227 9364 29239 9367
rect 29730 9364 29736 9376
rect 29227 9336 29736 9364
rect 29227 9333 29239 9336
rect 29181 9327 29239 9333
rect 29730 9324 29736 9336
rect 29788 9324 29794 9376
rect 31570 9324 31576 9376
rect 31628 9324 31634 9376
rect 31662 9324 31668 9376
rect 31720 9364 31726 9376
rect 33226 9364 33232 9376
rect 31720 9336 33232 9364
rect 31720 9324 31726 9336
rect 33226 9324 33232 9336
rect 33284 9324 33290 9376
rect 1104 9274 38272 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38272 9274
rect 1104 9200 38272 9222
rect 2958 9160 2964 9172
rect 2746 9132 2964 9160
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 2746 8956 2774 9132
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 6181 9163 6239 9169
rect 6181 9129 6193 9163
rect 6227 9160 6239 9163
rect 6822 9160 6828 9172
rect 6227 9132 6828 9160
rect 6227 9129 6239 9132
rect 6181 9123 6239 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 11517 9163 11575 9169
rect 7156 9132 11468 9160
rect 7156 9120 7162 9132
rect 3970 9052 3976 9104
rect 4028 9092 4034 9104
rect 6730 9092 6736 9104
rect 4028 9064 6736 9092
rect 4028 9052 4034 9064
rect 1811 8928 2774 8956
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 3326 8916 3332 8968
rect 3384 8916 3390 8968
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4264 8965 4292 9064
rect 6730 9052 6736 9064
rect 6788 9052 6794 9104
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 4356 8996 4629 9024
rect 4356 8965 4384 8996
rect 4617 8993 4629 8996
rect 4663 8993 4675 9027
rect 4617 8987 4675 8993
rect 4706 8984 4712 9036
rect 4764 9024 4770 9036
rect 7116 9024 7144 9120
rect 11440 9092 11468 9132
rect 11517 9129 11529 9163
rect 11563 9160 11575 9163
rect 11606 9160 11612 9172
rect 11563 9132 11612 9160
rect 11563 9129 11575 9132
rect 11517 9123 11575 9129
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 14090 9160 14096 9172
rect 12084 9132 14096 9160
rect 12084 9092 12112 9132
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 15286 9120 15292 9172
rect 15344 9160 15350 9172
rect 17497 9163 17555 9169
rect 17497 9160 17509 9163
rect 15344 9132 17509 9160
rect 15344 9120 15350 9132
rect 17497 9129 17509 9132
rect 17543 9160 17555 9163
rect 18230 9160 18236 9172
rect 17543 9132 18236 9160
rect 17543 9129 17555 9132
rect 17497 9123 17555 9129
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 18322 9120 18328 9172
rect 18380 9160 18386 9172
rect 19058 9160 19064 9172
rect 18380 9132 19064 9160
rect 18380 9120 18386 9132
rect 19058 9120 19064 9132
rect 19116 9120 19122 9172
rect 20901 9163 20959 9169
rect 20901 9129 20913 9163
rect 20947 9160 20959 9163
rect 21082 9160 21088 9172
rect 20947 9132 21088 9160
rect 20947 9129 20959 9132
rect 20901 9123 20959 9129
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 23937 9163 23995 9169
rect 23937 9160 23949 9163
rect 22152 9132 23949 9160
rect 22152 9120 22158 9132
rect 23937 9129 23949 9132
rect 23983 9160 23995 9163
rect 23983 9132 26188 9160
rect 23983 9129 23995 9132
rect 23937 9123 23995 9129
rect 11440 9064 12112 9092
rect 4764 8996 7144 9024
rect 8665 9027 8723 9033
rect 4764 8984 4770 8996
rect 8665 8993 8677 9027
rect 8711 9024 8723 9027
rect 9769 9027 9827 9033
rect 8711 8996 8800 9024
rect 8711 8993 8723 8996
rect 8665 8987 8723 8993
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8925 4399 8959
rect 4341 8919 4399 8925
rect 4525 8959 4583 8965
rect 4525 8925 4537 8959
rect 4571 8956 4583 8959
rect 4724 8956 4752 8984
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4571 8928 4752 8956
rect 4908 8928 4997 8956
rect 4571 8925 4583 8928
rect 4525 8919 4583 8925
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1397 8891 1455 8897
rect 1397 8888 1409 8891
rect 992 8860 1409 8888
rect 992 8848 998 8860
rect 1397 8857 1409 8860
rect 1443 8857 1455 8891
rect 3344 8888 3372 8916
rect 3344 8860 4660 8888
rect 1397 8851 1455 8857
rect 3878 8780 3884 8832
rect 3936 8780 3942 8832
rect 4632 8820 4660 8860
rect 4706 8848 4712 8900
rect 4764 8888 4770 8900
rect 4801 8891 4859 8897
rect 4801 8888 4813 8891
rect 4764 8860 4813 8888
rect 4764 8848 4770 8860
rect 4801 8857 4813 8860
rect 4847 8857 4859 8891
rect 4801 8851 4859 8857
rect 4908 8820 4936 8928
rect 4985 8925 4997 8928
rect 5031 8956 5043 8959
rect 5813 8959 5871 8965
rect 5813 8956 5825 8959
rect 5031 8928 5825 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5813 8925 5825 8928
rect 5859 8956 5871 8959
rect 7190 8956 7196 8968
rect 5859 8928 7196 8956
rect 5859 8925 5871 8928
rect 5813 8919 5871 8925
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 5994 8848 6000 8900
rect 6052 8848 6058 8900
rect 6178 8888 6184 8900
rect 6104 8860 6184 8888
rect 4632 8792 4936 8820
rect 5810 8780 5816 8832
rect 5868 8820 5874 8832
rect 6104 8820 6132 8860
rect 6178 8848 6184 8860
rect 6236 8888 6242 8900
rect 8772 8888 8800 8996
rect 9769 8993 9781 9027
rect 9815 8993 9827 9027
rect 9769 8987 9827 8993
rect 6236 8860 8800 8888
rect 9784 8888 9812 8987
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 10594 8984 10600 9036
rect 10652 9024 10658 9036
rect 13633 9027 13691 9033
rect 10652 8996 13492 9024
rect 10652 8984 10658 8996
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 12912 8965 12940 8996
rect 12713 8959 12771 8965
rect 12713 8956 12725 8959
rect 11388 8928 12725 8956
rect 11388 8916 11394 8928
rect 12713 8925 12725 8928
rect 12759 8925 12771 8959
rect 12713 8919 12771 8925
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8925 12955 8959
rect 12897 8919 12955 8925
rect 13354 8916 13360 8968
rect 13412 8916 13418 8968
rect 13464 8956 13492 8996
rect 13633 8993 13645 9027
rect 13679 9024 13691 9027
rect 13722 9024 13728 9036
rect 13679 8996 13728 9024
rect 13679 8993 13691 8996
rect 13633 8987 13691 8993
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 13814 8956 13820 8968
rect 13464 8928 13820 8956
rect 13814 8916 13820 8928
rect 13872 8916 13878 8968
rect 14108 8965 14136 9120
rect 14081 8959 14139 8965
rect 14081 8925 14093 8959
rect 14127 8925 14139 8959
rect 14081 8919 14139 8925
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 9950 8888 9956 8900
rect 9784 8860 9956 8888
rect 6236 8848 6242 8860
rect 5868 8792 6132 8820
rect 5868 8780 5874 8792
rect 8018 8780 8024 8832
rect 8076 8780 8082 8832
rect 8386 8780 8392 8832
rect 8444 8780 8450 8832
rect 8478 8780 8484 8832
rect 8536 8780 8542 8832
rect 8772 8820 8800 8860
rect 9950 8848 9956 8860
rect 10008 8848 10014 8900
rect 11422 8888 11428 8900
rect 11270 8860 11428 8888
rect 11422 8848 11428 8860
rect 11480 8848 11486 8900
rect 11698 8848 11704 8900
rect 11756 8848 11762 8900
rect 12805 8891 12863 8897
rect 12805 8857 12817 8891
rect 12851 8888 12863 8891
rect 14292 8888 14320 8919
rect 14366 8916 14372 8968
rect 14424 8956 14430 8968
rect 14507 8959 14565 8965
rect 14424 8928 14469 8956
rect 14424 8916 14430 8928
rect 14507 8925 14519 8959
rect 14553 8956 14565 8959
rect 15010 8956 15016 8968
rect 14553 8928 15016 8956
rect 14553 8925 14565 8928
rect 14507 8919 14565 8925
rect 15010 8916 15016 8928
rect 15068 8916 15074 8968
rect 15304 8965 15332 9120
rect 18966 9052 18972 9104
rect 19024 9092 19030 9104
rect 22833 9095 22891 9101
rect 19024 9064 22692 9092
rect 19024 9052 19030 9064
rect 15378 8984 15384 9036
rect 15436 9024 15442 9036
rect 15565 9027 15623 9033
rect 15565 9024 15577 9027
rect 15436 8996 15577 9024
rect 15436 8984 15442 8996
rect 15565 8993 15577 8996
rect 15611 9024 15623 9027
rect 17586 9024 17592 9036
rect 15611 8996 17592 9024
rect 15611 8993 15623 8996
rect 15565 8987 15623 8993
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 18325 9027 18383 9033
rect 18325 8993 18337 9027
rect 18371 8993 18383 9027
rect 20254 9024 20260 9036
rect 18325 8987 18383 8993
rect 19720 8996 20260 9024
rect 15289 8959 15347 8965
rect 15289 8925 15301 8959
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 15746 8916 15752 8968
rect 15804 8916 15810 8968
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 17328 8928 17969 8956
rect 12851 8860 14320 8888
rect 15381 8891 15439 8897
rect 12851 8857 12863 8860
rect 12805 8851 12863 8857
rect 15381 8857 15393 8891
rect 15427 8888 15439 8891
rect 15930 8888 15936 8900
rect 15427 8860 15936 8888
rect 15427 8857 15439 8860
rect 15381 8851 15439 8857
rect 15930 8848 15936 8860
rect 15988 8848 15994 8900
rect 16022 8848 16028 8900
rect 16080 8848 16086 8900
rect 16758 8848 16764 8900
rect 16816 8848 16822 8900
rect 11716 8820 11744 8848
rect 8772 8792 11744 8820
rect 12989 8823 13047 8829
rect 12989 8789 13001 8823
rect 13035 8820 13047 8823
rect 13078 8820 13084 8832
rect 13035 8792 13084 8820
rect 13035 8789 13047 8792
rect 12989 8783 13047 8789
rect 13078 8780 13084 8792
rect 13136 8780 13142 8832
rect 13446 8780 13452 8832
rect 13504 8820 13510 8832
rect 14642 8820 14648 8832
rect 13504 8792 14648 8820
rect 13504 8780 13510 8792
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 14734 8780 14740 8832
rect 14792 8780 14798 8832
rect 14918 8780 14924 8832
rect 14976 8780 14982 8832
rect 15948 8820 15976 8848
rect 17328 8820 17356 8928
rect 17957 8925 17969 8928
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 15948 8792 17356 8820
rect 18340 8820 18368 8987
rect 18690 8916 18696 8968
rect 18748 8916 18754 8968
rect 19720 8965 19748 8996
rect 20254 8984 20260 8996
rect 20312 8984 20318 9036
rect 20346 8984 20352 9036
rect 20404 9024 20410 9036
rect 20717 9027 20775 9033
rect 20717 9024 20729 9027
rect 20404 8996 20729 9024
rect 20404 8984 20410 8996
rect 20717 8993 20729 8996
rect 20763 8993 20775 9027
rect 20717 8987 20775 8993
rect 22186 8984 22192 9036
rect 22244 8984 22250 9036
rect 22664 9033 22692 9064
rect 22833 9061 22845 9095
rect 22879 9061 22891 9095
rect 22833 9055 22891 9061
rect 22649 9027 22707 9033
rect 22649 8993 22661 9027
rect 22695 8993 22707 9027
rect 22649 8987 22707 8993
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 19886 8916 19892 8968
rect 19944 8916 19950 8968
rect 19978 8916 19984 8968
rect 20036 8956 20042 8968
rect 20364 8956 20392 8984
rect 20036 8928 20392 8956
rect 20036 8916 20042 8928
rect 20622 8916 20628 8968
rect 20680 8916 20686 8968
rect 22554 8916 22560 8968
rect 22612 8916 22618 8968
rect 19521 8891 19579 8897
rect 19521 8857 19533 8891
rect 19567 8888 19579 8891
rect 20070 8888 20076 8900
rect 19567 8860 20076 8888
rect 19567 8857 19579 8860
rect 19521 8851 19579 8857
rect 20070 8848 20076 8860
rect 20128 8848 20134 8900
rect 20162 8848 20168 8900
rect 20220 8888 20226 8900
rect 20640 8888 20668 8916
rect 20220 8860 20668 8888
rect 20220 8848 20226 8860
rect 22278 8848 22284 8900
rect 22336 8848 22342 8900
rect 22664 8888 22692 8987
rect 22848 8956 22876 9055
rect 22922 9052 22928 9104
rect 22980 9052 22986 9104
rect 23106 9052 23112 9104
rect 23164 9092 23170 9104
rect 24394 9092 24400 9104
rect 23164 9064 24400 9092
rect 23164 9052 23170 9064
rect 24394 9052 24400 9064
rect 24452 9052 24458 9104
rect 24578 9052 24584 9104
rect 24636 9092 24642 9104
rect 24636 9064 24808 9092
rect 24636 9052 24642 9064
rect 22940 9024 22968 9052
rect 24780 9024 24808 9064
rect 24854 9052 24860 9104
rect 24912 9092 24918 9104
rect 26160 9092 26188 9132
rect 26602 9120 26608 9172
rect 26660 9160 26666 9172
rect 27246 9160 27252 9172
rect 26660 9132 27252 9160
rect 26660 9120 26666 9132
rect 27246 9120 27252 9132
rect 27304 9120 27310 9172
rect 29730 9120 29736 9172
rect 29788 9160 29794 9172
rect 29788 9132 30512 9160
rect 29788 9120 29794 9132
rect 27154 9092 27160 9104
rect 24912 9064 25636 9092
rect 24912 9052 24918 9064
rect 25317 9027 25375 9033
rect 22940 8996 24716 9024
rect 22925 8959 22983 8965
rect 22925 8956 22937 8959
rect 22848 8928 22937 8956
rect 22925 8925 22937 8928
rect 22971 8925 22983 8959
rect 22925 8919 22983 8925
rect 23014 8916 23020 8968
rect 23072 8956 23078 8968
rect 23216 8965 23244 8996
rect 23201 8959 23259 8965
rect 23072 8928 23117 8956
rect 23072 8916 23078 8928
rect 23201 8925 23213 8959
rect 23247 8925 23259 8959
rect 23201 8919 23259 8925
rect 23382 8916 23388 8968
rect 23440 8965 23446 8968
rect 23440 8956 23448 8965
rect 23440 8928 23485 8956
rect 23440 8919 23448 8928
rect 23440 8916 23446 8919
rect 23750 8916 23756 8968
rect 23808 8956 23814 8968
rect 23845 8959 23903 8965
rect 23845 8956 23857 8959
rect 23808 8928 23857 8956
rect 23808 8916 23814 8928
rect 23845 8925 23857 8928
rect 23891 8925 23903 8959
rect 23845 8919 23903 8925
rect 24394 8916 24400 8968
rect 24452 8916 24458 8968
rect 24688 8965 24716 8996
rect 24780 8996 25268 9024
rect 24780 8965 24808 8996
rect 24946 8965 24952 8968
rect 24490 8959 24548 8965
rect 24490 8925 24502 8959
rect 24536 8925 24548 8959
rect 24490 8919 24548 8925
rect 24673 8959 24731 8965
rect 24673 8925 24685 8959
rect 24719 8925 24731 8959
rect 24673 8919 24731 8925
rect 24765 8959 24823 8965
rect 24765 8925 24777 8959
rect 24811 8925 24823 8959
rect 24765 8919 24823 8925
rect 24903 8959 24952 8965
rect 24903 8925 24915 8959
rect 24949 8925 24952 8959
rect 24903 8919 24952 8925
rect 23290 8888 23296 8900
rect 22664 8860 23296 8888
rect 23290 8848 23296 8860
rect 23348 8888 23354 8900
rect 24504 8888 24532 8919
rect 24946 8916 24952 8919
rect 25004 8916 25010 8968
rect 25240 8965 25268 8996
rect 25317 8993 25329 9027
rect 25363 8993 25375 9027
rect 25317 8987 25375 8993
rect 25225 8959 25283 8965
rect 25225 8925 25237 8959
rect 25271 8925 25283 8959
rect 25225 8919 25283 8925
rect 24578 8888 24584 8900
rect 23348 8860 24584 8888
rect 23348 8848 23354 8860
rect 24578 8848 24584 8860
rect 24636 8848 24642 8900
rect 20346 8820 20352 8832
rect 18340 8792 20352 8820
rect 20346 8780 20352 8792
rect 20404 8820 20410 8832
rect 21818 8820 21824 8832
rect 20404 8792 21824 8820
rect 20404 8780 20410 8792
rect 21818 8780 21824 8792
rect 21876 8780 21882 8832
rect 23566 8780 23572 8832
rect 23624 8780 23630 8832
rect 25041 8823 25099 8829
rect 25041 8789 25053 8823
rect 25087 8820 25099 8823
rect 25130 8820 25136 8832
rect 25087 8792 25136 8820
rect 25087 8789 25099 8792
rect 25041 8783 25099 8789
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 25240 8820 25268 8919
rect 25332 8900 25360 8987
rect 25406 8916 25412 8968
rect 25464 8956 25470 8968
rect 25608 8965 25636 9064
rect 26160 9064 27160 9092
rect 25777 9027 25835 9033
rect 25777 8993 25789 9027
rect 25823 9024 25835 9027
rect 25823 8996 26096 9024
rect 25823 8993 25835 8996
rect 25777 8987 25835 8993
rect 25501 8959 25559 8965
rect 25501 8956 25513 8959
rect 25464 8928 25513 8956
rect 25464 8916 25470 8928
rect 25501 8925 25513 8928
rect 25547 8925 25559 8959
rect 25501 8919 25559 8925
rect 25593 8959 25651 8965
rect 25593 8925 25605 8959
rect 25639 8925 25651 8959
rect 25593 8919 25651 8925
rect 25866 8916 25872 8968
rect 25924 8916 25930 8968
rect 26068 8965 26096 8996
rect 26160 8965 26188 9064
rect 27154 9052 27160 9064
rect 27212 9052 27218 9104
rect 29178 9092 29184 9104
rect 27816 9064 29184 9092
rect 27816 9036 27844 9064
rect 26510 9024 26516 9036
rect 26252 8996 26516 9024
rect 26252 8965 26280 8996
rect 26510 8984 26516 8996
rect 26568 9024 26574 9036
rect 27065 9027 27123 9033
rect 27065 9024 27077 9027
rect 26568 8996 26740 9024
rect 26568 8984 26574 8996
rect 26053 8959 26111 8965
rect 26053 8925 26065 8959
rect 26099 8925 26111 8959
rect 26053 8919 26111 8925
rect 26145 8959 26203 8965
rect 26145 8925 26157 8959
rect 26191 8925 26203 8959
rect 26145 8919 26203 8925
rect 26237 8959 26295 8965
rect 26237 8925 26249 8959
rect 26283 8925 26295 8959
rect 26237 8919 26295 8925
rect 25314 8848 25320 8900
rect 25372 8888 25378 8900
rect 25774 8888 25780 8900
rect 25372 8860 25780 8888
rect 25372 8848 25378 8860
rect 25774 8848 25780 8860
rect 25832 8888 25838 8900
rect 26712 8888 26740 8996
rect 26896 8996 27077 9024
rect 26786 8916 26792 8968
rect 26844 8916 26850 8968
rect 26896 8888 26924 8996
rect 27065 8993 27077 8996
rect 27111 8993 27123 9027
rect 27065 8987 27123 8993
rect 27798 8984 27804 9036
rect 27856 8984 27862 9036
rect 28074 8984 28080 9036
rect 28132 8984 28138 9036
rect 26970 8916 26976 8968
rect 27028 8916 27034 8968
rect 27154 8916 27160 8968
rect 27212 8916 27218 8968
rect 27246 8916 27252 8968
rect 27304 8956 27310 8968
rect 27341 8959 27399 8965
rect 27341 8956 27353 8959
rect 27304 8928 27353 8956
rect 27304 8916 27310 8928
rect 27341 8925 27353 8928
rect 27387 8925 27399 8959
rect 27341 8919 27399 8925
rect 27617 8959 27675 8965
rect 27617 8925 27629 8959
rect 27663 8925 27675 8959
rect 27617 8919 27675 8925
rect 27632 8888 27660 8919
rect 27982 8916 27988 8968
rect 28040 8916 28046 8968
rect 28092 8956 28120 8984
rect 28169 8959 28227 8965
rect 28169 8956 28181 8959
rect 28092 8928 28181 8956
rect 28169 8925 28181 8928
rect 28215 8925 28227 8959
rect 28169 8919 28227 8925
rect 28353 8959 28411 8965
rect 28353 8925 28365 8959
rect 28399 8925 28411 8959
rect 28353 8919 28411 8925
rect 25832 8860 26648 8888
rect 26712 8860 26924 8888
rect 26988 8860 27660 8888
rect 25832 8848 25838 8860
rect 26326 8820 26332 8832
rect 25240 8792 26332 8820
rect 26326 8780 26332 8792
rect 26384 8780 26390 8832
rect 26510 8780 26516 8832
rect 26568 8780 26574 8832
rect 26620 8820 26648 8860
rect 26988 8820 27016 8860
rect 27706 8848 27712 8900
rect 27764 8888 27770 8900
rect 27801 8891 27859 8897
rect 27801 8888 27813 8891
rect 27764 8860 27813 8888
rect 27764 8848 27770 8860
rect 27801 8857 27813 8860
rect 27847 8857 27859 8891
rect 28368 8888 28396 8919
rect 28442 8916 28448 8968
rect 28500 8916 28506 8968
rect 28920 8965 28948 9064
rect 29178 9052 29184 9064
rect 29236 9052 29242 9104
rect 29822 9052 29828 9104
rect 29880 9052 29886 9104
rect 29917 9095 29975 9101
rect 29917 9061 29929 9095
rect 29963 9061 29975 9095
rect 29917 9055 29975 9061
rect 29273 9027 29331 9033
rect 29012 8996 29224 9024
rect 28537 8959 28595 8965
rect 28537 8925 28549 8959
rect 28583 8925 28595 8959
rect 28537 8919 28595 8925
rect 28905 8959 28963 8965
rect 28905 8925 28917 8959
rect 28951 8925 28963 8959
rect 28905 8919 28963 8925
rect 27801 8851 27859 8857
rect 27908 8860 28396 8888
rect 28552 8888 28580 8919
rect 28552 8860 28948 8888
rect 26620 8792 27016 8820
rect 27525 8823 27583 8829
rect 27525 8789 27537 8823
rect 27571 8820 27583 8823
rect 27908 8820 27936 8860
rect 28920 8832 28948 8860
rect 29012 8832 29040 8996
rect 29196 8965 29224 8996
rect 29273 8993 29285 9027
rect 29319 9024 29331 9027
rect 29840 9024 29868 9052
rect 29319 8996 29868 9024
rect 29319 8993 29331 8996
rect 29273 8987 29331 8993
rect 29089 8959 29147 8965
rect 29089 8925 29101 8959
rect 29135 8925 29147 8959
rect 29089 8919 29147 8925
rect 29187 8959 29245 8965
rect 29187 8925 29199 8959
rect 29233 8925 29245 8959
rect 29187 8919 29245 8925
rect 29104 8888 29132 8919
rect 29362 8916 29368 8968
rect 29420 8916 29426 8968
rect 29564 8965 29592 8996
rect 29549 8959 29607 8965
rect 29549 8925 29561 8959
rect 29595 8925 29607 8959
rect 29549 8919 29607 8925
rect 29641 8959 29699 8965
rect 29641 8925 29653 8959
rect 29687 8925 29699 8959
rect 29932 8956 29960 9055
rect 30009 8959 30067 8965
rect 30009 8956 30021 8959
rect 29932 8928 30021 8956
rect 29641 8919 29699 8925
rect 30009 8925 30021 8928
rect 30055 8925 30067 8959
rect 30009 8919 30067 8925
rect 29270 8888 29276 8900
rect 29104 8860 29276 8888
rect 29270 8848 29276 8860
rect 29328 8848 29334 8900
rect 27571 8792 27936 8820
rect 27571 8789 27583 8792
rect 27525 8783 27583 8789
rect 28810 8780 28816 8832
rect 28868 8780 28874 8832
rect 28902 8780 28908 8832
rect 28960 8780 28966 8832
rect 28994 8780 29000 8832
rect 29052 8780 29058 8832
rect 29086 8780 29092 8832
rect 29144 8820 29150 8832
rect 29656 8820 29684 8919
rect 30098 8916 30104 8968
rect 30156 8956 30162 8968
rect 30193 8959 30251 8965
rect 30193 8956 30205 8959
rect 30156 8928 30205 8956
rect 30156 8916 30162 8928
rect 30193 8925 30205 8928
rect 30239 8925 30251 8959
rect 30193 8919 30251 8925
rect 30374 8848 30380 8900
rect 30432 8848 30438 8900
rect 30484 8888 30512 9132
rect 30742 9120 30748 9172
rect 30800 9120 30806 9172
rect 31570 9120 31576 9172
rect 31628 9160 31634 9172
rect 31757 9163 31815 9169
rect 31757 9160 31769 9163
rect 31628 9132 31769 9160
rect 31628 9120 31634 9132
rect 31757 9129 31769 9132
rect 31803 9129 31815 9163
rect 31757 9123 31815 9129
rect 32861 9163 32919 9169
rect 32861 9129 32873 9163
rect 32907 9160 32919 9163
rect 33134 9160 33140 9172
rect 32907 9132 33140 9160
rect 32907 9129 32919 9132
rect 32861 9123 32919 9129
rect 33134 9120 33140 9132
rect 33192 9120 33198 9172
rect 33229 9163 33287 9169
rect 33229 9129 33241 9163
rect 33275 9160 33287 9163
rect 33318 9160 33324 9172
rect 33275 9132 33324 9160
rect 33275 9129 33287 9132
rect 33229 9123 33287 9129
rect 33318 9120 33324 9132
rect 33376 9120 33382 9172
rect 30760 9092 30788 9120
rect 32401 9095 32459 9101
rect 32401 9092 32413 9095
rect 30760 9064 32413 9092
rect 32401 9061 32413 9064
rect 32447 9061 32459 9095
rect 32401 9055 32459 9061
rect 32784 9064 33548 9092
rect 31481 9027 31539 9033
rect 31481 8993 31493 9027
rect 31527 9024 31539 9027
rect 32030 9024 32036 9036
rect 31527 8996 32036 9024
rect 31527 8993 31539 8996
rect 31481 8987 31539 8993
rect 32030 8984 32036 8996
rect 32088 8984 32094 9036
rect 32784 8968 32812 9064
rect 33520 9033 33548 9064
rect 33505 9027 33563 9033
rect 33505 8993 33517 9027
rect 33551 8993 33563 9027
rect 33505 8987 33563 8993
rect 31573 8959 31631 8965
rect 31573 8925 31585 8959
rect 31619 8956 31631 8959
rect 31754 8956 31760 8968
rect 31619 8928 31760 8956
rect 31619 8925 31631 8928
rect 31573 8919 31631 8925
rect 31754 8916 31760 8928
rect 31812 8916 31818 8968
rect 31846 8916 31852 8968
rect 31904 8916 31910 8968
rect 32125 8959 32183 8965
rect 32125 8925 32137 8959
rect 32171 8956 32183 8959
rect 32585 8959 32643 8965
rect 32171 8928 32536 8956
rect 32171 8925 32183 8928
rect 32125 8919 32183 8925
rect 32140 8888 32168 8919
rect 30484 8860 32168 8888
rect 29144 8792 29684 8820
rect 29144 8780 29150 8792
rect 30926 8780 30932 8832
rect 30984 8820 30990 8832
rect 31113 8823 31171 8829
rect 31113 8820 31125 8823
rect 30984 8792 31125 8820
rect 30984 8780 30990 8792
rect 31113 8789 31125 8792
rect 31159 8789 31171 8823
rect 31113 8783 31171 8789
rect 31938 8780 31944 8832
rect 31996 8780 32002 8832
rect 32508 8820 32536 8928
rect 32585 8925 32597 8959
rect 32631 8925 32643 8959
rect 32585 8919 32643 8925
rect 32677 8959 32735 8965
rect 32677 8925 32689 8959
rect 32723 8956 32735 8959
rect 32766 8956 32772 8968
rect 32723 8928 32772 8956
rect 32723 8925 32735 8928
rect 32677 8919 32735 8925
rect 32600 8888 32628 8919
rect 32766 8916 32772 8928
rect 32824 8916 32830 8968
rect 32953 8959 33011 8965
rect 32953 8925 32965 8959
rect 32999 8925 33011 8959
rect 32953 8919 33011 8925
rect 32858 8888 32864 8900
rect 32600 8860 32864 8888
rect 32858 8848 32864 8860
rect 32916 8848 32922 8900
rect 32968 8888 32996 8919
rect 33042 8916 33048 8968
rect 33100 8916 33106 8968
rect 33134 8916 33140 8968
rect 33192 8916 33198 8968
rect 33229 8959 33287 8965
rect 33229 8925 33241 8959
rect 33275 8925 33287 8959
rect 33229 8919 33287 8925
rect 37921 8959 37979 8965
rect 37921 8925 37933 8959
rect 37967 8956 37979 8959
rect 38286 8956 38292 8968
rect 37967 8928 38292 8956
rect 37967 8925 37979 8928
rect 37921 8919 37979 8925
rect 33152 8888 33180 8916
rect 32968 8860 33180 8888
rect 33244 8832 33272 8919
rect 38286 8916 38292 8928
rect 38344 8916 38350 8968
rect 35894 8848 35900 8900
rect 35952 8888 35958 8900
rect 36814 8888 36820 8900
rect 35952 8860 36820 8888
rect 35952 8848 35958 8860
rect 36814 8848 36820 8860
rect 36872 8888 36878 8900
rect 37645 8891 37703 8897
rect 37645 8888 37657 8891
rect 36872 8860 37657 8888
rect 36872 8848 36878 8860
rect 37645 8857 37657 8860
rect 37691 8857 37703 8891
rect 37645 8851 37703 8857
rect 33226 8820 33232 8832
rect 32508 8792 33232 8820
rect 33226 8780 33232 8792
rect 33284 8780 33290 8832
rect 1104 8730 38272 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38272 8730
rect 1104 8656 38272 8678
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 4295 8588 5089 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 5077 8579 5135 8585
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 6365 8619 6423 8625
rect 6365 8616 6377 8619
rect 5960 8588 6377 8616
rect 5960 8576 5966 8588
rect 6365 8585 6377 8588
rect 6411 8585 6423 8619
rect 6365 8579 6423 8585
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 9677 8619 9735 8625
rect 9677 8616 9689 8619
rect 8536 8588 9689 8616
rect 8536 8576 8542 8588
rect 9677 8585 9689 8588
rect 9723 8585 9735 8619
rect 9677 8579 9735 8585
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 10134 8616 10140 8628
rect 10091 8588 10140 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 10428 8588 10609 8616
rect 6517 8551 6575 8557
rect 6517 8548 6529 8551
rect 4724 8520 6529 8548
rect 4724 8492 4752 8520
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8480 3479 8483
rect 4157 8483 4215 8489
rect 3467 8452 3832 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 3804 8353 3832 8452
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4706 8480 4712 8492
rect 4203 8452 4712 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 5920 8489 5948 8520
rect 6517 8517 6529 8520
rect 6563 8517 6575 8551
rect 6517 8511 6575 8517
rect 6733 8551 6791 8557
rect 6733 8517 6745 8551
rect 6779 8517 6791 8551
rect 6733 8511 6791 8517
rect 7837 8551 7895 8557
rect 7837 8517 7849 8551
rect 7883 8548 7895 8551
rect 7883 8520 9996 8548
rect 7883 8517 7895 8520
rect 7837 8511 7895 8517
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4479 8384 4752 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 3789 8347 3847 8353
rect 3789 8313 3801 8347
rect 3835 8313 3847 8347
rect 3789 8307 3847 8313
rect 4062 8304 4068 8356
rect 4120 8344 4126 8356
rect 4120 8316 4660 8344
rect 4120 8304 4126 8316
rect 4632 8288 4660 8316
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3237 8279 3295 8285
rect 3237 8276 3249 8279
rect 3016 8248 3249 8276
rect 3016 8236 3022 8248
rect 3237 8245 3249 8248
rect 3283 8245 3295 8279
rect 3237 8239 3295 8245
rect 4614 8236 4620 8288
rect 4672 8236 4678 8288
rect 4724 8276 4752 8384
rect 5460 8344 5488 8443
rect 5994 8440 6000 8492
rect 6052 8480 6058 8492
rect 6089 8483 6147 8489
rect 6089 8480 6101 8483
rect 6052 8452 6101 8480
rect 6052 8440 6058 8452
rect 6089 8449 6101 8452
rect 6135 8449 6147 8483
rect 6089 8443 6147 8449
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8480 6239 8483
rect 6362 8480 6368 8492
rect 6227 8452 6368 8480
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 5534 8372 5540 8424
rect 5592 8372 5598 8424
rect 5626 8372 5632 8424
rect 5684 8372 5690 8424
rect 6104 8412 6132 8443
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 6748 8412 6776 8511
rect 9968 8492 9996 8520
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 9585 8483 9643 8489
rect 9585 8480 9597 8483
rect 9456 8452 9597 8480
rect 9456 8440 9462 8452
rect 9585 8449 9597 8452
rect 9631 8480 9643 8483
rect 9858 8480 9864 8492
rect 9631 8452 9864 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 9858 8440 9864 8452
rect 9916 8440 9922 8492
rect 9950 8440 9956 8492
rect 10008 8440 10014 8492
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8480 10195 8483
rect 10428 8480 10456 8588
rect 10597 8585 10609 8588
rect 10643 8616 10655 8619
rect 11330 8616 11336 8628
rect 10643 8588 11336 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 12250 8576 12256 8628
rect 12308 8616 12314 8628
rect 12308 8588 13492 8616
rect 12308 8576 12314 8588
rect 12437 8551 12495 8557
rect 12437 8548 12449 8551
rect 11992 8520 12449 8548
rect 10183 8452 10456 8480
rect 10183 8449 10195 8452
rect 10137 8443 10195 8449
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11204 8452 11529 8480
rect 11204 8440 11210 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 11992 8489 12020 8520
rect 12437 8517 12449 8520
rect 12483 8517 12495 8551
rect 12437 8511 12495 8517
rect 12618 8508 12624 8560
rect 12676 8508 12682 8560
rect 13078 8508 13084 8560
rect 13136 8508 13142 8560
rect 11977 8483 12035 8489
rect 11977 8480 11989 8483
rect 11848 8452 11989 8480
rect 11848 8440 11854 8452
rect 11977 8449 11989 8452
rect 12023 8449 12035 8483
rect 11977 8443 12035 8449
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8449 12403 8483
rect 12345 8443 12403 8449
rect 6104 8384 6776 8412
rect 10321 8415 10379 8421
rect 10321 8381 10333 8415
rect 10367 8412 10379 8415
rect 10410 8412 10416 8424
rect 10367 8384 10416 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 11882 8372 11888 8424
rect 11940 8372 11946 8424
rect 12158 8344 12164 8356
rect 5460 8316 12164 8344
rect 12158 8304 12164 8316
rect 12216 8304 12222 8356
rect 5718 8276 5724 8288
rect 4724 8248 5724 8276
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 5902 8236 5908 8288
rect 5960 8236 5966 8288
rect 6362 8236 6368 8288
rect 6420 8276 6426 8288
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 6420 8248 6561 8276
rect 6420 8236 6426 8248
rect 6549 8245 6561 8248
rect 6595 8276 6607 8279
rect 6822 8276 6828 8288
rect 6595 8248 6828 8276
rect 6595 8245 6607 8248
rect 6549 8239 6607 8245
rect 6822 8236 6828 8248
rect 6880 8276 6886 8288
rect 8386 8276 8392 8288
rect 6880 8248 8392 8276
rect 6880 8236 6886 8248
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 12360 8276 12388 8443
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 13096 8480 13124 8508
rect 13464 8489 13492 8588
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 15197 8619 15255 8625
rect 15197 8616 15209 8619
rect 14700 8588 15209 8616
rect 14700 8576 14706 8588
rect 15197 8585 15209 8588
rect 15243 8616 15255 8619
rect 18414 8616 18420 8628
rect 15243 8588 18420 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 18877 8619 18935 8625
rect 18877 8585 18889 8619
rect 18923 8616 18935 8619
rect 18966 8616 18972 8628
rect 18923 8588 18972 8616
rect 18923 8585 18935 8588
rect 18877 8579 18935 8585
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 20254 8616 20260 8628
rect 19536 8588 20260 8616
rect 17310 8508 17316 8560
rect 17368 8548 17374 8560
rect 19536 8557 19564 8588
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 21818 8576 21824 8628
rect 21876 8616 21882 8628
rect 21876 8588 23152 8616
rect 21876 8576 21882 8588
rect 19521 8551 19579 8557
rect 17368 8520 19472 8548
rect 17368 8508 17374 8520
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 13096 8452 13185 8480
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 13173 8443 13231 8449
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8449 13507 8483
rect 16758 8480 16764 8492
rect 14858 8452 16764 8480
rect 13449 8443 13507 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17494 8440 17500 8492
rect 17552 8440 17558 8492
rect 18598 8440 18604 8492
rect 18656 8480 18662 8492
rect 18785 8483 18843 8489
rect 18785 8480 18797 8483
rect 18656 8452 18797 8480
rect 18656 8440 18662 8452
rect 18785 8449 18797 8452
rect 18831 8480 18843 8483
rect 18874 8480 18880 8492
rect 18831 8452 18880 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 18966 8440 18972 8492
rect 19024 8440 19030 8492
rect 19444 8480 19472 8520
rect 19521 8517 19533 8551
rect 19567 8517 19579 8551
rect 19521 8511 19579 8517
rect 19628 8520 21588 8548
rect 19628 8480 19656 8520
rect 19444 8452 19656 8480
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8449 19763 8483
rect 19705 8443 19763 8449
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8480 19855 8483
rect 19978 8480 19984 8492
rect 19843 8452 19984 8480
rect 19843 8449 19855 8452
rect 19797 8443 19855 8449
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 13372 8384 13737 8412
rect 13372 8353 13400 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 15010 8372 15016 8424
rect 15068 8412 15074 8424
rect 19720 8412 19748 8443
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 20162 8412 20168 8424
rect 15068 8384 19334 8412
rect 19720 8384 20168 8412
rect 15068 8372 15074 8384
rect 13357 8347 13415 8353
rect 13357 8313 13369 8347
rect 13403 8313 13415 8347
rect 13357 8307 13415 8313
rect 17218 8304 17224 8356
rect 17276 8304 17282 8356
rect 19306 8344 19334 8384
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 21560 8412 21588 8520
rect 21634 8508 21640 8560
rect 21692 8548 21698 8560
rect 22097 8551 22155 8557
rect 22097 8548 22109 8551
rect 21692 8520 22109 8548
rect 21692 8508 21698 8520
rect 22097 8517 22109 8520
rect 22143 8517 22155 8551
rect 22097 8511 22155 8517
rect 21913 8483 21971 8489
rect 21913 8449 21925 8483
rect 21959 8480 21971 8483
rect 22002 8480 22008 8492
rect 21959 8452 22008 8480
rect 21959 8449 21971 8452
rect 21913 8443 21971 8449
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 23124 8412 23152 8588
rect 23566 8576 23572 8628
rect 23624 8576 23630 8628
rect 24302 8576 24308 8628
rect 24360 8616 24366 8628
rect 24949 8619 25007 8625
rect 24949 8616 24961 8619
rect 24360 8588 24961 8616
rect 24360 8576 24366 8588
rect 24949 8585 24961 8588
rect 24995 8616 25007 8619
rect 26970 8616 26976 8628
rect 24995 8588 26976 8616
rect 24995 8585 25007 8588
rect 24949 8579 25007 8585
rect 26970 8576 26976 8588
rect 27028 8576 27034 8628
rect 28902 8576 28908 8628
rect 28960 8616 28966 8628
rect 29273 8619 29331 8625
rect 28960 8588 29132 8616
rect 28960 8576 28966 8588
rect 23584 8548 23612 8576
rect 23216 8520 23612 8548
rect 23216 8489 23244 8520
rect 24118 8508 24124 8560
rect 24176 8548 24182 8560
rect 24176 8520 24900 8548
rect 24176 8508 24182 8520
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8449 23259 8483
rect 23201 8443 23259 8449
rect 23477 8483 23535 8489
rect 23477 8449 23489 8483
rect 23523 8480 23535 8483
rect 23566 8480 23572 8492
rect 23523 8452 23572 8480
rect 23523 8449 23535 8452
rect 23477 8443 23535 8449
rect 23566 8440 23572 8452
rect 23624 8440 23630 8492
rect 23661 8483 23719 8489
rect 23661 8449 23673 8483
rect 23707 8480 23719 8483
rect 23842 8480 23848 8492
rect 23707 8452 23848 8480
rect 23707 8449 23719 8452
rect 23661 8443 23719 8449
rect 23842 8440 23848 8452
rect 23900 8480 23906 8492
rect 24670 8480 24676 8492
rect 23900 8452 24676 8480
rect 23900 8440 23906 8452
rect 24670 8440 24676 8452
rect 24728 8440 24734 8492
rect 24872 8489 24900 8520
rect 25314 8508 25320 8560
rect 25372 8508 25378 8560
rect 26988 8548 27016 8576
rect 28994 8548 29000 8560
rect 26988 8520 27200 8548
rect 24857 8483 24915 8489
rect 24857 8449 24869 8483
rect 24903 8480 24915 8483
rect 25332 8480 25360 8508
rect 24903 8452 25360 8480
rect 24903 8449 24915 8452
rect 24857 8443 24915 8449
rect 26510 8440 26516 8492
rect 26568 8480 26574 8492
rect 27172 8489 27200 8520
rect 27264 8520 29000 8548
rect 27264 8489 27292 8520
rect 28994 8508 29000 8520
rect 29052 8508 29058 8560
rect 29104 8548 29132 8588
rect 29273 8585 29285 8619
rect 29319 8616 29331 8619
rect 30098 8616 30104 8628
rect 29319 8588 30104 8616
rect 29319 8585 29331 8588
rect 29273 8579 29331 8585
rect 30098 8576 30104 8588
rect 30156 8576 30162 8628
rect 31297 8619 31355 8625
rect 31297 8585 31309 8619
rect 31343 8616 31355 8619
rect 31386 8616 31392 8628
rect 31343 8588 31392 8616
rect 31343 8585 31355 8588
rect 31297 8579 31355 8585
rect 31386 8576 31392 8588
rect 31444 8576 31450 8628
rect 32030 8576 32036 8628
rect 32088 8576 32094 8628
rect 30190 8548 30196 8560
rect 29104 8520 30196 8548
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26568 8452 26985 8480
rect 26568 8440 26574 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27157 8483 27215 8489
rect 27157 8449 27169 8483
rect 27203 8449 27215 8483
rect 27157 8443 27215 8449
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8449 27307 8483
rect 27249 8443 27307 8449
rect 27341 8483 27399 8489
rect 27341 8449 27353 8483
rect 27387 8449 27399 8483
rect 27341 8443 27399 8449
rect 27525 8483 27583 8489
rect 27525 8449 27537 8483
rect 27571 8449 27583 8483
rect 27525 8443 27583 8449
rect 23290 8412 23296 8424
rect 21560 8384 22094 8412
rect 23124 8384 23296 8412
rect 21910 8344 21916 8356
rect 19306 8316 21916 8344
rect 21910 8304 21916 8316
rect 21968 8304 21974 8356
rect 22066 8344 22094 8384
rect 23290 8372 23296 8384
rect 23348 8412 23354 8424
rect 24765 8415 24823 8421
rect 24765 8412 24777 8415
rect 23348 8384 24777 8412
rect 23348 8372 23354 8384
rect 24765 8381 24777 8384
rect 24811 8412 24823 8415
rect 25406 8412 25412 8424
rect 24811 8384 25412 8412
rect 24811 8381 24823 8384
rect 24765 8375 24823 8381
rect 25406 8372 25412 8384
rect 25464 8372 25470 8424
rect 26786 8372 26792 8424
rect 26844 8412 26850 8424
rect 27062 8412 27068 8424
rect 26844 8384 27068 8412
rect 26844 8372 26850 8384
rect 27062 8372 27068 8384
rect 27120 8412 27126 8424
rect 27356 8412 27384 8443
rect 27120 8384 27384 8412
rect 27120 8372 27126 8384
rect 27540 8356 27568 8443
rect 27614 8440 27620 8492
rect 27672 8480 27678 8492
rect 29104 8489 29132 8520
rect 30190 8508 30196 8520
rect 30248 8548 30254 8560
rect 31938 8548 31944 8560
rect 30248 8520 31944 8548
rect 30248 8508 30254 8520
rect 31938 8508 31944 8520
rect 31996 8508 32002 8560
rect 28905 8483 28963 8489
rect 28905 8480 28917 8483
rect 27672 8452 28917 8480
rect 27672 8440 27678 8452
rect 28905 8449 28917 8452
rect 28951 8449 28963 8483
rect 28905 8443 28963 8449
rect 29089 8483 29147 8489
rect 29089 8449 29101 8483
rect 29135 8449 29147 8483
rect 29089 8443 29147 8449
rect 31573 8483 31631 8489
rect 31573 8449 31585 8483
rect 31619 8480 31631 8483
rect 31662 8480 31668 8492
rect 31619 8452 31668 8480
rect 31619 8449 31631 8452
rect 31573 8443 31631 8449
rect 28920 8412 28948 8443
rect 31662 8440 31668 8452
rect 31720 8440 31726 8492
rect 31849 8483 31907 8489
rect 31849 8449 31861 8483
rect 31895 8480 31907 8483
rect 32048 8480 32076 8576
rect 35894 8548 35900 8560
rect 31895 8452 32076 8480
rect 32968 8520 35900 8548
rect 31895 8449 31907 8452
rect 31849 8443 31907 8449
rect 29362 8412 29368 8424
rect 28920 8384 29368 8412
rect 29362 8372 29368 8384
rect 29420 8372 29426 8424
rect 31018 8372 31024 8424
rect 31076 8412 31082 8424
rect 31389 8415 31447 8421
rect 31389 8412 31401 8415
rect 31076 8384 31401 8412
rect 31076 8372 31082 8384
rect 31389 8381 31401 8384
rect 31435 8381 31447 8415
rect 32968 8412 32996 8520
rect 35894 8508 35900 8520
rect 35952 8508 35958 8560
rect 33042 8440 33048 8492
rect 33100 8480 33106 8492
rect 33137 8483 33195 8489
rect 33137 8480 33149 8483
rect 33100 8452 33149 8480
rect 33100 8440 33106 8452
rect 33137 8449 33149 8452
rect 33183 8449 33195 8483
rect 33137 8443 33195 8449
rect 31389 8375 31447 8381
rect 31726 8384 32996 8412
rect 22066 8316 27476 8344
rect 12802 8276 12808 8288
rect 12360 8248 12808 8276
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 13722 8236 13728 8288
rect 13780 8276 13786 8288
rect 15654 8276 15660 8288
rect 13780 8248 15660 8276
rect 13780 8236 13786 8248
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 19518 8236 19524 8288
rect 19576 8236 19582 8288
rect 22281 8279 22339 8285
rect 22281 8245 22293 8279
rect 22327 8276 22339 8279
rect 22370 8276 22376 8288
rect 22327 8248 22376 8276
rect 22327 8245 22339 8248
rect 22281 8239 22339 8245
rect 22370 8236 22376 8248
rect 22428 8236 22434 8288
rect 23014 8236 23020 8288
rect 23072 8236 23078 8288
rect 25314 8236 25320 8288
rect 25372 8236 25378 8288
rect 27448 8276 27476 8316
rect 27522 8304 27528 8356
rect 27580 8304 27586 8356
rect 27709 8347 27767 8353
rect 27709 8313 27721 8347
rect 27755 8344 27767 8347
rect 27798 8344 27804 8356
rect 27755 8316 27804 8344
rect 27755 8313 27767 8316
rect 27709 8307 27767 8313
rect 27798 8304 27804 8316
rect 27856 8304 27862 8356
rect 31726 8344 31754 8384
rect 33226 8372 33232 8424
rect 33284 8372 33290 8424
rect 27908 8316 31754 8344
rect 27908 8276 27936 8316
rect 32582 8304 32588 8356
rect 32640 8344 32646 8356
rect 32769 8347 32827 8353
rect 32769 8344 32781 8347
rect 32640 8316 32781 8344
rect 32640 8304 32646 8316
rect 32769 8313 32781 8316
rect 32815 8313 32827 8347
rect 32769 8307 32827 8313
rect 27448 8248 27936 8276
rect 28994 8236 29000 8288
rect 29052 8236 29058 8288
rect 29638 8236 29644 8288
rect 29696 8276 29702 8288
rect 34054 8276 34060 8288
rect 29696 8248 34060 8276
rect 29696 8236 29702 8248
rect 34054 8236 34060 8248
rect 34112 8236 34118 8288
rect 1104 8186 38272 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38272 8186
rect 1104 8112 38272 8134
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 5629 8075 5687 8081
rect 5629 8072 5641 8075
rect 5592 8044 5641 8072
rect 5592 8032 5598 8044
rect 5629 8041 5641 8044
rect 5675 8041 5687 8075
rect 5629 8035 5687 8041
rect 5810 8032 5816 8084
rect 5868 8032 5874 8084
rect 6472 8044 8248 8072
rect 5828 7936 5856 8032
rect 5644 7908 5856 7936
rect 5644 7877 5672 7908
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5718 7828 5724 7880
rect 5776 7828 5782 7880
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7868 5871 7871
rect 5902 7868 5908 7880
rect 5859 7840 5908 7868
rect 5859 7837 5871 7840
rect 5813 7831 5871 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6472 7877 6500 8044
rect 8220 8004 8248 8044
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 8665 8075 8723 8081
rect 8665 8072 8677 8075
rect 8444 8044 8677 8072
rect 8444 8032 8450 8044
rect 8665 8041 8677 8044
rect 8711 8072 8723 8075
rect 10502 8072 10508 8084
rect 8711 8044 10508 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 11885 8075 11943 8081
rect 11885 8072 11897 8075
rect 11572 8044 11897 8072
rect 11572 8032 11578 8044
rect 11885 8041 11897 8044
rect 11931 8072 11943 8075
rect 12250 8072 12256 8084
rect 11931 8044 12256 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 12805 8075 12863 8081
rect 12805 8072 12817 8075
rect 12584 8044 12817 8072
rect 12584 8032 12590 8044
rect 12805 8041 12817 8044
rect 12851 8041 12863 8075
rect 12805 8035 12863 8041
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 13541 8075 13599 8081
rect 13541 8072 13553 8075
rect 13044 8044 13553 8072
rect 13044 8032 13050 8044
rect 13541 8041 13553 8044
rect 13587 8041 13599 8075
rect 13541 8035 13599 8041
rect 13722 8032 13728 8084
rect 13780 8032 13786 8084
rect 19426 8032 19432 8084
rect 19484 8032 19490 8084
rect 20165 8075 20223 8081
rect 20165 8041 20177 8075
rect 20211 8072 20223 8075
rect 23566 8072 23572 8084
rect 20211 8044 23572 8072
rect 20211 8041 20223 8044
rect 20165 8035 20223 8041
rect 23566 8032 23572 8044
rect 23624 8032 23630 8084
rect 26234 8032 26240 8084
rect 26292 8072 26298 8084
rect 29270 8072 29276 8084
rect 26292 8044 29276 8072
rect 26292 8032 26298 8044
rect 29270 8032 29276 8044
rect 29328 8032 29334 8084
rect 30834 8032 30840 8084
rect 30892 8072 30898 8084
rect 31478 8072 31484 8084
rect 30892 8044 31484 8072
rect 30892 8032 30898 8044
rect 31478 8032 31484 8044
rect 31536 8032 31542 8084
rect 31754 8032 31760 8084
rect 31812 8072 31818 8084
rect 31849 8075 31907 8081
rect 31849 8072 31861 8075
rect 31812 8044 31861 8072
rect 31812 8032 31818 8044
rect 31849 8041 31861 8044
rect 31895 8041 31907 8075
rect 31849 8035 31907 8041
rect 17497 8007 17555 8013
rect 17497 8004 17509 8007
rect 8220 7976 17509 8004
rect 17497 7973 17509 7976
rect 17543 7973 17555 8007
rect 19444 8004 19472 8032
rect 20254 8004 20260 8016
rect 19444 7976 20260 8004
rect 17497 7967 17555 7973
rect 20254 7964 20260 7976
rect 20312 7964 20318 8016
rect 21637 8007 21695 8013
rect 21637 7973 21649 8007
rect 21683 8004 21695 8007
rect 22646 8004 22652 8016
rect 21683 7976 22652 8004
rect 21683 7973 21695 7976
rect 21637 7967 21695 7973
rect 22646 7964 22652 7976
rect 22704 7964 22710 8016
rect 22738 7964 22744 8016
rect 22796 8004 22802 8016
rect 23293 8007 23351 8013
rect 23293 8004 23305 8007
rect 22796 7976 23305 8004
rect 22796 7964 22802 7976
rect 23293 7973 23305 7976
rect 23339 7973 23351 8007
rect 23293 7967 23351 7973
rect 24026 7964 24032 8016
rect 24084 8004 24090 8016
rect 30745 8007 30803 8013
rect 24084 7976 30604 8004
rect 24084 7964 24090 7976
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 5736 7800 5764 7828
rect 6656 7800 6684 7899
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 9398 7936 9404 7948
rect 6972 7908 9404 7936
rect 6972 7896 6978 7908
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 11882 7936 11888 7948
rect 9784 7908 11888 7936
rect 9674 7828 9680 7880
rect 9732 7877 9738 7880
rect 9732 7868 9743 7877
rect 9784 7868 9812 7908
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 12621 7939 12679 7945
rect 12621 7905 12633 7939
rect 12667 7936 12679 7939
rect 13630 7936 13636 7948
rect 12667 7908 13636 7936
rect 12667 7905 12679 7908
rect 12621 7899 12679 7905
rect 9732 7840 9812 7868
rect 9861 7871 9919 7877
rect 9732 7831 9743 7840
rect 9861 7837 9873 7871
rect 9907 7837 9919 7871
rect 9861 7831 9919 7837
rect 9732 7828 9738 7831
rect 5736 7772 6684 7800
rect 7190 7760 7196 7812
rect 7248 7760 7254 7812
rect 8478 7800 8484 7812
rect 8418 7772 8484 7800
rect 8478 7760 8484 7772
rect 8536 7800 8542 7812
rect 9766 7800 9772 7812
rect 8536 7772 9772 7800
rect 8536 7760 8542 7772
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 6086 7692 6092 7744
rect 6144 7692 6150 7744
rect 6546 7692 6552 7744
rect 6604 7692 6610 7744
rect 9674 7692 9680 7744
rect 9732 7692 9738 7744
rect 9876 7732 9904 7831
rect 9950 7828 9956 7880
rect 10008 7868 10014 7880
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 10008 7840 10425 7868
rect 10008 7828 10014 7840
rect 10413 7837 10425 7840
rect 10459 7868 10471 7871
rect 10962 7868 10968 7880
rect 10459 7840 10968 7868
rect 10459 7837 10471 7840
rect 10413 7831 10471 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 12342 7760 12348 7812
rect 12400 7760 12406 7812
rect 10870 7732 10876 7744
rect 9876 7704 10876 7732
rect 10870 7692 10876 7704
rect 10928 7732 10934 7744
rect 12636 7732 12664 7899
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 13998 7896 14004 7948
rect 14056 7896 14062 7948
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 15933 7939 15991 7945
rect 15933 7936 15945 7939
rect 15712 7908 15945 7936
rect 15712 7896 15718 7908
rect 15933 7905 15945 7908
rect 15979 7905 15991 7939
rect 15933 7899 15991 7905
rect 17144 7908 17816 7936
rect 13354 7828 13360 7880
rect 13412 7868 13418 7880
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13412 7840 13737 7868
rect 13412 7828 13418 7840
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7837 13967 7871
rect 14016 7868 14044 7896
rect 15749 7871 15807 7877
rect 15749 7868 15761 7871
rect 14016 7840 15761 7868
rect 13909 7831 13967 7837
rect 15749 7837 15761 7840
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7868 15899 7871
rect 17144 7868 17172 7908
rect 17788 7880 17816 7908
rect 19518 7896 19524 7948
rect 19576 7896 19582 7948
rect 20622 7936 20628 7948
rect 19904 7908 20628 7936
rect 15887 7840 17172 7868
rect 17221 7871 17279 7877
rect 15887 7837 15899 7840
rect 15841 7831 15899 7837
rect 17221 7837 17233 7871
rect 17267 7868 17279 7871
rect 17586 7868 17592 7880
rect 17267 7840 17592 7868
rect 17267 7837 17279 7840
rect 17221 7831 17279 7837
rect 13630 7760 13636 7812
rect 13688 7800 13694 7812
rect 13924 7800 13952 7831
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 17770 7828 17776 7880
rect 17828 7828 17834 7880
rect 19536 7868 19564 7896
rect 19904 7877 19932 7908
rect 20622 7896 20628 7908
rect 20680 7936 20686 7948
rect 22278 7936 22284 7948
rect 20680 7908 22284 7936
rect 20680 7896 20686 7908
rect 19705 7871 19763 7877
rect 19705 7868 19717 7871
rect 19536 7840 19717 7868
rect 19705 7837 19717 7840
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 19889 7871 19947 7877
rect 19889 7837 19901 7871
rect 19935 7837 19947 7871
rect 19889 7831 19947 7837
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7868 20315 7871
rect 21545 7871 21603 7877
rect 20303 7840 20576 7868
rect 20303 7837 20315 7840
rect 20257 7831 20315 7837
rect 16850 7800 16856 7812
rect 13688 7772 16856 7800
rect 13688 7760 13694 7772
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 17497 7803 17555 7809
rect 17497 7769 17509 7803
rect 17543 7800 17555 7803
rect 17681 7803 17739 7809
rect 17681 7800 17693 7803
rect 17543 7772 17693 7800
rect 17543 7769 17555 7772
rect 17497 7763 17555 7769
rect 17681 7769 17693 7772
rect 17727 7769 17739 7803
rect 17681 7763 17739 7769
rect 19797 7803 19855 7809
rect 19797 7769 19809 7803
rect 19843 7800 19855 7803
rect 20088 7800 20116 7831
rect 19843 7772 20116 7800
rect 19843 7769 19855 7772
rect 19797 7763 19855 7769
rect 20548 7744 20576 7840
rect 21545 7837 21557 7871
rect 21591 7868 21603 7871
rect 21634 7868 21640 7880
rect 21591 7840 21640 7868
rect 21591 7837 21603 7840
rect 21545 7831 21603 7837
rect 21634 7828 21640 7840
rect 21692 7828 21698 7880
rect 21744 7877 21772 7908
rect 22278 7896 22284 7908
rect 22336 7896 22342 7948
rect 22370 7896 22376 7948
rect 22428 7896 22434 7948
rect 23014 7936 23020 7948
rect 22572 7908 23020 7936
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7837 21787 7871
rect 21729 7831 21787 7837
rect 21818 7828 21824 7880
rect 21876 7828 21882 7880
rect 21913 7871 21971 7877
rect 21913 7837 21925 7871
rect 21959 7837 21971 7871
rect 21913 7831 21971 7837
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7837 22155 7871
rect 22097 7831 22155 7837
rect 22189 7871 22247 7877
rect 22189 7837 22201 7871
rect 22235 7868 22247 7871
rect 22572 7868 22600 7908
rect 23014 7896 23020 7908
rect 23072 7896 23078 7948
rect 28994 7896 29000 7948
rect 29052 7936 29058 7948
rect 29914 7936 29920 7948
rect 29052 7908 29920 7936
rect 29052 7896 29058 7908
rect 29914 7896 29920 7908
rect 29972 7936 29978 7948
rect 30285 7939 30343 7945
rect 29972 7908 30236 7936
rect 29972 7896 29978 7908
rect 22235 7840 22600 7868
rect 22235 7837 22247 7840
rect 22189 7831 22247 7837
rect 10928 7704 12664 7732
rect 10928 7692 10934 7704
rect 15378 7692 15384 7744
rect 15436 7692 15442 7744
rect 17310 7692 17316 7744
rect 17368 7692 17374 7744
rect 20530 7692 20536 7744
rect 20588 7692 20594 7744
rect 21928 7732 21956 7831
rect 22112 7800 22140 7831
rect 22646 7828 22652 7880
rect 22704 7828 22710 7880
rect 30006 7828 30012 7880
rect 30064 7828 30070 7880
rect 30208 7877 30236 7908
rect 30285 7905 30297 7939
rect 30331 7936 30343 7939
rect 30466 7936 30472 7948
rect 30331 7908 30472 7936
rect 30331 7905 30343 7908
rect 30285 7899 30343 7905
rect 30466 7896 30472 7908
rect 30524 7896 30530 7948
rect 30576 7936 30604 7976
rect 30745 7973 30757 8007
rect 30791 8004 30803 8007
rect 33042 8004 33048 8016
rect 30791 7976 33048 8004
rect 30791 7973 30803 7976
rect 30745 7967 30803 7973
rect 33042 7964 33048 7976
rect 33100 7964 33106 8016
rect 31110 7936 31116 7948
rect 30576 7908 31116 7936
rect 31110 7896 31116 7908
rect 31168 7896 31174 7948
rect 30193 7871 30251 7877
rect 30193 7837 30205 7871
rect 30239 7837 30251 7871
rect 30193 7831 30251 7837
rect 30374 7828 30380 7880
rect 30432 7828 30438 7880
rect 30561 7871 30619 7877
rect 30561 7868 30573 7871
rect 30484 7840 30573 7868
rect 22370 7800 22376 7812
rect 22112 7772 22376 7800
rect 22370 7760 22376 7772
rect 22428 7760 22434 7812
rect 22554 7760 22560 7812
rect 22612 7800 22618 7812
rect 22741 7803 22799 7809
rect 22741 7800 22753 7803
rect 22612 7772 22753 7800
rect 22612 7760 22618 7772
rect 22741 7769 22753 7772
rect 22787 7769 22799 7803
rect 22741 7763 22799 7769
rect 23106 7760 23112 7812
rect 23164 7760 23170 7812
rect 25038 7760 25044 7812
rect 25096 7800 25102 7812
rect 25866 7800 25872 7812
rect 25096 7772 25872 7800
rect 25096 7760 25102 7772
rect 25866 7760 25872 7772
rect 25924 7800 25930 7812
rect 27338 7800 27344 7812
rect 25924 7772 27344 7800
rect 25924 7760 25930 7772
rect 27338 7760 27344 7772
rect 27396 7800 27402 7812
rect 30484 7800 30512 7840
rect 30561 7837 30573 7840
rect 30607 7868 30619 7871
rect 30834 7868 30840 7880
rect 30607 7840 30840 7868
rect 30607 7837 30619 7840
rect 30561 7831 30619 7837
rect 30834 7828 30840 7840
rect 30892 7828 30898 7880
rect 30926 7828 30932 7880
rect 30984 7828 30990 7880
rect 31018 7828 31024 7880
rect 31076 7868 31082 7880
rect 31389 7871 31447 7877
rect 31389 7868 31401 7871
rect 31076 7840 31401 7868
rect 31076 7828 31082 7840
rect 31389 7837 31401 7840
rect 31435 7868 31447 7871
rect 31481 7871 31539 7877
rect 31481 7868 31493 7871
rect 31435 7840 31493 7868
rect 31435 7837 31447 7840
rect 31389 7831 31447 7837
rect 31481 7837 31493 7840
rect 31527 7837 31539 7871
rect 31481 7831 31539 7837
rect 31297 7803 31355 7809
rect 31297 7800 31309 7803
rect 27396 7772 30512 7800
rect 30576 7772 31309 7800
rect 27396 7760 27402 7772
rect 30576 7744 30604 7772
rect 31297 7769 31309 7772
rect 31343 7800 31355 7803
rect 31662 7800 31668 7812
rect 31343 7772 31668 7800
rect 31343 7769 31355 7772
rect 31297 7763 31355 7769
rect 31662 7760 31668 7772
rect 31720 7760 31726 7812
rect 22094 7732 22100 7744
rect 21928 7704 22100 7732
rect 22094 7692 22100 7704
rect 22152 7692 22158 7744
rect 22278 7692 22284 7744
rect 22336 7692 22342 7744
rect 30558 7692 30564 7744
rect 30616 7692 30622 7744
rect 31202 7692 31208 7744
rect 31260 7692 31266 7744
rect 1104 7642 38272 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38272 7642
rect 1104 7568 38272 7590
rect 4614 7528 4620 7540
rect 2608 7500 4620 7528
rect 1486 7352 1492 7404
rect 1544 7352 1550 7404
rect 2608 7401 2636 7500
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 5629 7531 5687 7537
rect 5629 7497 5641 7531
rect 5675 7528 5687 7531
rect 6086 7528 6092 7540
rect 5675 7500 6092 7528
rect 5675 7497 5687 7500
rect 5629 7491 5687 7497
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 6546 7488 6552 7540
rect 6604 7488 6610 7540
rect 7190 7488 7196 7540
rect 7248 7528 7254 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 7248 7500 7665 7528
rect 7248 7488 7254 7500
rect 7653 7497 7665 7500
rect 7699 7497 7711 7531
rect 7653 7491 7711 7497
rect 8018 7488 8024 7540
rect 8076 7488 8082 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13228 7500 14872 7528
rect 13228 7488 13234 7500
rect 2869 7463 2927 7469
rect 2869 7429 2881 7463
rect 2915 7460 2927 7463
rect 2958 7460 2964 7472
rect 2915 7432 2964 7460
rect 2915 7429 2927 7432
rect 2869 7423 2927 7429
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 3970 7352 3976 7404
rect 4028 7352 4034 7404
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7392 5595 7395
rect 5994 7392 6000 7404
rect 5583 7364 6000 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 3602 7324 3608 7336
rect 1719 7296 3608 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 4341 7327 4399 7333
rect 4341 7293 4353 7327
rect 4387 7324 4399 7327
rect 4706 7324 4712 7336
rect 4387 7296 4712 7324
rect 4387 7293 4399 7296
rect 4341 7287 4399 7293
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7293 5871 7327
rect 5813 7287 5871 7293
rect 5166 7148 5172 7200
rect 5224 7148 5230 7200
rect 5828 7188 5856 7287
rect 6012 7256 6040 7352
rect 6365 7327 6423 7333
rect 6365 7293 6377 7327
rect 6411 7324 6423 7327
rect 6564 7324 6592 7488
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8036 7392 8064 7488
rect 9766 7420 9772 7472
rect 9824 7460 9830 7472
rect 9824 7432 10166 7460
rect 9824 7420 9830 7432
rect 11790 7420 11796 7472
rect 11848 7420 11854 7472
rect 12434 7420 12440 7472
rect 12492 7420 12498 7472
rect 14642 7460 14648 7472
rect 14568 7432 14648 7460
rect 14568 7401 14596 7432
rect 14642 7420 14648 7432
rect 14700 7420 14706 7472
rect 14844 7401 14872 7500
rect 15378 7488 15384 7540
rect 15436 7488 15442 7540
rect 18598 7488 18604 7540
rect 18656 7488 18662 7540
rect 19613 7531 19671 7537
rect 19613 7528 19625 7531
rect 18708 7500 19625 7528
rect 7883 7364 8064 7392
rect 14553 7395 14611 7401
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 14553 7361 14565 7395
rect 14599 7361 14611 7395
rect 14553 7355 14611 7361
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7392 14887 7395
rect 15286 7392 15292 7404
rect 14875 7364 15292 7392
rect 14875 7361 14887 7364
rect 14829 7355 14887 7361
rect 6411 7296 6592 7324
rect 6411 7293 6423 7296
rect 6365 7287 6423 7293
rect 6748 7256 6776 7355
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15396 7392 15424 7488
rect 18616 7460 18644 7488
rect 18708 7472 18736 7500
rect 19613 7497 19625 7500
rect 19659 7528 19671 7531
rect 21358 7528 21364 7540
rect 19659 7500 21364 7528
rect 19659 7497 19671 7500
rect 19613 7491 19671 7497
rect 21358 7488 21364 7500
rect 21416 7488 21422 7540
rect 22278 7488 22284 7540
rect 22336 7488 22342 7540
rect 22370 7488 22376 7540
rect 22428 7488 22434 7540
rect 22756 7500 23060 7528
rect 17972 7432 18644 7460
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15396 7364 15485 7392
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 17770 7352 17776 7404
rect 17828 7352 17834 7404
rect 17972 7401 18000 7432
rect 18690 7420 18696 7472
rect 18748 7420 18754 7472
rect 19337 7463 19395 7469
rect 19337 7429 19349 7463
rect 19383 7460 19395 7463
rect 20165 7463 20223 7469
rect 20165 7460 20177 7463
rect 19383 7432 20177 7460
rect 19383 7429 19395 7432
rect 19337 7423 19395 7429
rect 20165 7429 20177 7432
rect 20211 7429 20223 7463
rect 20165 7423 20223 7429
rect 17957 7395 18015 7401
rect 17957 7361 17969 7395
rect 18003 7361 18015 7395
rect 19153 7395 19211 7401
rect 19153 7392 19165 7395
rect 17957 7355 18015 7361
rect 18064 7364 19165 7392
rect 6822 7284 6828 7336
rect 6880 7284 6886 7336
rect 9398 7284 9404 7336
rect 9456 7284 9462 7336
rect 9674 7284 9680 7336
rect 9732 7284 9738 7336
rect 11514 7284 11520 7336
rect 11572 7284 11578 7336
rect 14274 7284 14280 7336
rect 14332 7324 14338 7336
rect 14461 7327 14519 7333
rect 14461 7324 14473 7327
rect 14332 7296 14473 7324
rect 14332 7284 14338 7296
rect 14461 7293 14473 7296
rect 14507 7324 14519 7327
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 14507 7296 14657 7324
rect 14507 7293 14519 7296
rect 14461 7287 14519 7293
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 15013 7327 15071 7333
rect 15013 7293 15025 7327
rect 15059 7324 15071 7327
rect 15378 7324 15384 7336
rect 15059 7296 15384 7324
rect 15059 7293 15071 7296
rect 15013 7287 15071 7293
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 6012 7228 6776 7256
rect 13538 7216 13544 7268
rect 13596 7256 13602 7268
rect 14185 7259 14243 7265
rect 14185 7256 14197 7259
rect 13596 7228 14197 7256
rect 13596 7216 13602 7228
rect 14185 7225 14197 7228
rect 14231 7225 14243 7259
rect 14185 7219 14243 7225
rect 18064 7200 18092 7364
rect 19153 7361 19165 7364
rect 19199 7392 19211 7395
rect 19521 7395 19579 7401
rect 19521 7392 19533 7395
rect 19199 7364 19533 7392
rect 19199 7361 19211 7364
rect 19153 7355 19211 7361
rect 19521 7361 19533 7364
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 19797 7395 19855 7401
rect 19797 7361 19809 7395
rect 19843 7361 19855 7395
rect 19797 7355 19855 7361
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7392 20407 7395
rect 20622 7392 20628 7404
rect 20395 7364 20628 7392
rect 20395 7361 20407 7364
rect 20349 7355 20407 7361
rect 18690 7284 18696 7336
rect 18748 7324 18754 7336
rect 18969 7327 19027 7333
rect 18969 7324 18981 7327
rect 18748 7296 18981 7324
rect 18748 7284 18754 7296
rect 18969 7293 18981 7296
rect 19015 7293 19027 7327
rect 18969 7287 19027 7293
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 19812 7324 19840 7355
rect 20622 7352 20628 7364
rect 20680 7392 20686 7404
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 20680 7364 20821 7392
rect 20680 7352 20686 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 21376 7392 21404 7488
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 21376 7364 21833 7392
rect 20809 7355 20867 7361
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 22094 7352 22100 7404
rect 22152 7352 22158 7404
rect 22186 7352 22192 7404
rect 22244 7352 22250 7404
rect 22296 7392 22324 7488
rect 22756 7401 22784 7500
rect 22922 7420 22928 7472
rect 22980 7420 22986 7472
rect 23032 7460 23060 7500
rect 23106 7488 23112 7540
rect 23164 7528 23170 7540
rect 23201 7531 23259 7537
rect 23201 7528 23213 7531
rect 23164 7500 23213 7528
rect 23164 7488 23170 7500
rect 23201 7497 23213 7500
rect 23247 7497 23259 7531
rect 26418 7528 26424 7540
rect 23201 7491 23259 7497
rect 23860 7500 26424 7528
rect 23860 7460 23888 7500
rect 26418 7488 26424 7500
rect 26476 7488 26482 7540
rect 26602 7488 26608 7540
rect 26660 7528 26666 7540
rect 27522 7528 27528 7540
rect 26660 7500 27528 7528
rect 26660 7488 26666 7500
rect 27522 7488 27528 7500
rect 27580 7488 27586 7540
rect 27614 7488 27620 7540
rect 27672 7488 27678 7540
rect 27706 7488 27712 7540
rect 27764 7528 27770 7540
rect 27764 7500 29500 7528
rect 27764 7488 27770 7500
rect 23032 7432 23888 7460
rect 23937 7463 23995 7469
rect 23937 7429 23949 7463
rect 23983 7460 23995 7463
rect 25038 7460 25044 7472
rect 23983 7432 24164 7460
rect 23983 7429 23995 7432
rect 23937 7423 23995 7429
rect 22557 7395 22615 7401
rect 22557 7392 22569 7395
rect 22296 7364 22569 7392
rect 22557 7361 22569 7364
rect 22603 7361 22615 7395
rect 22557 7355 22615 7361
rect 22705 7395 22784 7401
rect 22705 7361 22717 7395
rect 22751 7364 22784 7395
rect 22833 7395 22891 7401
rect 22751 7361 22763 7364
rect 22705 7355 22763 7361
rect 22833 7361 22845 7395
rect 22879 7361 22891 7395
rect 22833 7355 22891 7361
rect 23063 7395 23121 7401
rect 23063 7361 23075 7395
rect 23109 7392 23121 7395
rect 23109 7364 23244 7392
rect 23109 7361 23121 7364
rect 23063 7355 23121 7361
rect 19484 7296 19840 7324
rect 20901 7327 20959 7333
rect 19484 7284 19490 7296
rect 20901 7293 20913 7327
rect 20947 7324 20959 7327
rect 21082 7324 21088 7336
rect 20947 7296 21088 7324
rect 20947 7293 20959 7296
rect 20901 7287 20959 7293
rect 21082 7284 21088 7296
rect 21140 7284 21146 7336
rect 21266 7284 21272 7336
rect 21324 7324 21330 7336
rect 22848 7324 22876 7355
rect 21324 7296 22876 7324
rect 23216 7324 23244 7364
rect 23566 7352 23572 7404
rect 23624 7392 23630 7404
rect 23845 7395 23903 7401
rect 23845 7392 23857 7395
rect 23624 7364 23857 7392
rect 23624 7352 23630 7364
rect 23845 7361 23857 7364
rect 23891 7361 23903 7395
rect 23845 7355 23903 7361
rect 24026 7352 24032 7404
rect 24084 7352 24090 7404
rect 24136 7401 24164 7432
rect 24320 7432 25044 7460
rect 24320 7401 24348 7432
rect 25038 7420 25044 7432
rect 25096 7420 25102 7472
rect 25314 7420 25320 7472
rect 25372 7460 25378 7472
rect 25593 7463 25651 7469
rect 25593 7460 25605 7463
rect 25372 7432 25605 7460
rect 25372 7420 25378 7432
rect 25593 7429 25605 7432
rect 25639 7429 25651 7463
rect 25593 7423 25651 7429
rect 26234 7420 26240 7472
rect 26292 7420 26298 7472
rect 26326 7420 26332 7472
rect 26384 7460 26390 7472
rect 26384 7432 26648 7460
rect 26384 7420 26390 7432
rect 24121 7395 24179 7401
rect 24121 7361 24133 7395
rect 24167 7361 24179 7395
rect 24121 7355 24179 7361
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 24486 7352 24492 7404
rect 24544 7352 24550 7404
rect 24578 7352 24584 7404
rect 24636 7392 24642 7404
rect 24673 7395 24731 7401
rect 24673 7392 24685 7395
rect 24636 7364 24685 7392
rect 24636 7352 24642 7364
rect 24673 7361 24685 7364
rect 24719 7361 24731 7395
rect 24673 7355 24731 7361
rect 25133 7395 25191 7401
rect 25133 7361 25145 7395
rect 25179 7392 25191 7395
rect 25222 7392 25228 7404
rect 25179 7364 25228 7392
rect 25179 7361 25191 7364
rect 25133 7355 25191 7361
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 26252 7392 26280 7420
rect 26620 7401 26648 7432
rect 27338 7420 27344 7472
rect 27396 7420 27402 7472
rect 27632 7460 27660 7488
rect 27632 7432 27844 7460
rect 26421 7395 26479 7401
rect 26421 7392 26433 7395
rect 26252 7364 26433 7392
rect 26421 7361 26433 7364
rect 26467 7361 26479 7395
rect 26421 7355 26479 7361
rect 26605 7395 26663 7401
rect 26605 7361 26617 7395
rect 26651 7361 26663 7395
rect 27356 7392 27384 7420
rect 27816 7401 27844 7432
rect 27617 7395 27675 7401
rect 27617 7392 27629 7395
rect 27356 7364 27629 7392
rect 26605 7355 26663 7361
rect 27617 7361 27629 7364
rect 27663 7361 27675 7395
rect 27617 7355 27675 7361
rect 27801 7395 27859 7401
rect 27801 7361 27813 7395
rect 27847 7361 27859 7395
rect 27801 7355 27859 7361
rect 27893 7395 27951 7401
rect 27893 7361 27905 7395
rect 27939 7361 27951 7395
rect 27893 7355 27951 7361
rect 27985 7395 28043 7401
rect 27985 7361 27997 7395
rect 28031 7392 28043 7395
rect 28445 7395 28503 7401
rect 28445 7392 28457 7395
rect 28031 7364 28457 7392
rect 28031 7361 28043 7364
rect 27985 7355 28043 7361
rect 28445 7361 28457 7364
rect 28491 7392 28503 7395
rect 28534 7392 28540 7404
rect 28491 7364 28540 7392
rect 28491 7361 28503 7364
rect 28445 7355 28503 7361
rect 24397 7327 24455 7333
rect 24397 7324 24409 7327
rect 23216 7296 24409 7324
rect 21324 7284 21330 7296
rect 19981 7259 20039 7265
rect 19981 7225 19993 7259
rect 20027 7256 20039 7259
rect 21177 7259 21235 7265
rect 20027 7228 20576 7256
rect 20027 7225 20039 7228
rect 19981 7219 20039 7225
rect 20548 7200 20576 7228
rect 21177 7225 21189 7259
rect 21223 7256 21235 7259
rect 22002 7256 22008 7268
rect 21223 7228 22008 7256
rect 21223 7225 21235 7228
rect 21177 7219 21235 7225
rect 22002 7216 22008 7228
rect 22060 7256 22066 7268
rect 23216 7256 23244 7296
rect 24397 7293 24409 7296
rect 24443 7293 24455 7327
rect 24397 7287 24455 7293
rect 25317 7327 25375 7333
rect 25317 7293 25329 7327
rect 25363 7324 25375 7327
rect 25406 7324 25412 7336
rect 25363 7296 25412 7324
rect 25363 7293 25375 7296
rect 25317 7287 25375 7293
rect 25406 7284 25412 7296
rect 25464 7284 25470 7336
rect 27709 7327 27767 7333
rect 27709 7293 27721 7327
rect 27755 7324 27767 7327
rect 27908 7324 27936 7355
rect 28534 7352 28540 7364
rect 28592 7352 28598 7404
rect 28994 7352 29000 7404
rect 29052 7352 29058 7404
rect 29089 7395 29147 7401
rect 29089 7361 29101 7395
rect 29135 7361 29147 7395
rect 29089 7355 29147 7361
rect 27755 7296 27936 7324
rect 27755 7293 27767 7296
rect 27709 7287 27767 7293
rect 28258 7284 28264 7336
rect 28316 7284 28322 7336
rect 22060 7228 23244 7256
rect 22060 7216 22066 7228
rect 23566 7216 23572 7268
rect 23624 7256 23630 7268
rect 23624 7228 28028 7256
rect 23624 7216 23630 7228
rect 6178 7188 6184 7200
rect 5828 7160 6184 7188
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 11146 7148 11152 7200
rect 11204 7148 11210 7200
rect 12894 7148 12900 7200
rect 12952 7188 12958 7200
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 12952 7160 13277 7188
rect 12952 7148 12958 7160
rect 13265 7157 13277 7160
rect 13311 7188 13323 7191
rect 13354 7188 13360 7200
rect 13311 7160 13360 7188
rect 13311 7157 13323 7160
rect 13265 7151 13323 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 14553 7191 14611 7197
rect 14553 7157 14565 7191
rect 14599 7188 14611 7191
rect 14918 7188 14924 7200
rect 14599 7160 14924 7188
rect 14599 7157 14611 7160
rect 14553 7151 14611 7157
rect 14918 7148 14924 7160
rect 14976 7188 14982 7200
rect 15470 7188 15476 7200
rect 14976 7160 15476 7188
rect 14976 7148 14982 7160
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 15562 7148 15568 7200
rect 15620 7188 15626 7200
rect 15657 7191 15715 7197
rect 15657 7188 15669 7191
rect 15620 7160 15669 7188
rect 15620 7148 15626 7160
rect 15657 7157 15669 7160
rect 15703 7157 15715 7191
rect 15657 7151 15715 7157
rect 17862 7148 17868 7200
rect 17920 7148 17926 7200
rect 18046 7148 18052 7200
rect 18104 7148 18110 7200
rect 20530 7148 20536 7200
rect 20588 7148 20594 7200
rect 20898 7148 20904 7200
rect 20956 7188 20962 7200
rect 21913 7191 21971 7197
rect 21913 7188 21925 7191
rect 20956 7160 21925 7188
rect 20956 7148 20962 7160
rect 21913 7157 21925 7160
rect 21959 7188 21971 7191
rect 24486 7188 24492 7200
rect 21959 7160 24492 7188
rect 21959 7157 21971 7160
rect 21913 7151 21971 7157
rect 24486 7148 24492 7160
rect 24544 7148 24550 7200
rect 24854 7148 24860 7200
rect 24912 7148 24918 7200
rect 24949 7191 25007 7197
rect 24949 7157 24961 7191
rect 24995 7188 25007 7191
rect 25038 7188 25044 7200
rect 24995 7160 25044 7188
rect 24995 7157 25007 7160
rect 24949 7151 25007 7157
rect 25038 7148 25044 7160
rect 25096 7148 25102 7200
rect 25130 7148 25136 7200
rect 25188 7148 25194 7200
rect 26694 7148 26700 7200
rect 26752 7188 26758 7200
rect 27706 7188 27712 7200
rect 26752 7160 27712 7188
rect 26752 7148 26758 7160
rect 27706 7148 27712 7160
rect 27764 7148 27770 7200
rect 28000 7188 28028 7228
rect 28074 7216 28080 7268
rect 28132 7256 28138 7268
rect 29104 7256 29132 7355
rect 29178 7352 29184 7404
rect 29236 7392 29242 7404
rect 29365 7395 29423 7401
rect 29365 7392 29377 7395
rect 29236 7364 29377 7392
rect 29236 7352 29242 7364
rect 29365 7361 29377 7364
rect 29411 7361 29423 7395
rect 29365 7355 29423 7361
rect 29472 7324 29500 7500
rect 29638 7488 29644 7540
rect 29696 7488 29702 7540
rect 30006 7488 30012 7540
rect 30064 7528 30070 7540
rect 30101 7531 30159 7537
rect 30101 7528 30113 7531
rect 30064 7500 30113 7528
rect 30064 7488 30070 7500
rect 30101 7497 30113 7500
rect 30147 7497 30159 7531
rect 30101 7491 30159 7497
rect 31202 7488 31208 7540
rect 31260 7528 31266 7540
rect 31260 7500 31754 7528
rect 31260 7488 31266 7500
rect 29656 7401 29684 7488
rect 31570 7460 31576 7472
rect 30300 7432 31576 7460
rect 30300 7401 30328 7432
rect 31570 7420 31576 7432
rect 31628 7420 31634 7472
rect 31726 7460 31754 7500
rect 31726 7432 31892 7460
rect 29641 7395 29699 7401
rect 29641 7361 29653 7395
rect 29687 7361 29699 7395
rect 29641 7355 29699 7361
rect 30101 7395 30159 7401
rect 30101 7361 30113 7395
rect 30147 7361 30159 7395
rect 30285 7395 30343 7401
rect 30285 7392 30297 7395
rect 30101 7355 30159 7361
rect 30208 7364 30297 7392
rect 30116 7324 30144 7355
rect 29472 7296 30144 7324
rect 28132 7228 29132 7256
rect 28132 7216 28138 7228
rect 30208 7188 30236 7364
rect 30285 7361 30297 7364
rect 30331 7361 30343 7395
rect 30285 7355 30343 7361
rect 30650 7352 30656 7404
rect 30708 7392 30714 7404
rect 30745 7395 30803 7401
rect 30745 7392 30757 7395
rect 30708 7364 30757 7392
rect 30708 7352 30714 7364
rect 30745 7361 30757 7364
rect 30791 7361 30803 7395
rect 30745 7355 30803 7361
rect 31386 7352 31392 7404
rect 31444 7352 31450 7404
rect 31754 7352 31760 7404
rect 31812 7352 31818 7404
rect 31864 7401 31892 7432
rect 31849 7395 31907 7401
rect 31849 7361 31861 7395
rect 31895 7361 31907 7395
rect 31849 7355 31907 7361
rect 31294 7284 31300 7336
rect 31352 7284 31358 7336
rect 28000 7160 30236 7188
rect 1104 7098 38272 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38272 7098
rect 1104 7024 38272 7046
rect 5994 6944 6000 6996
rect 6052 6944 6058 6996
rect 12342 6944 12348 6996
rect 12400 6944 12406 6996
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 13630 6984 13636 6996
rect 12860 6956 13636 6984
rect 12860 6944 12866 6956
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 15562 6944 15568 6996
rect 15620 6984 15626 6996
rect 15730 6987 15788 6993
rect 15730 6984 15742 6987
rect 15620 6956 15742 6984
rect 15620 6944 15626 6956
rect 15730 6953 15742 6956
rect 15776 6953 15788 6987
rect 15730 6947 15788 6953
rect 17221 6987 17279 6993
rect 17221 6953 17233 6987
rect 17267 6984 17279 6987
rect 17770 6984 17776 6996
rect 17267 6956 17776 6984
rect 17267 6953 17279 6956
rect 17221 6947 17279 6953
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 18046 6944 18052 6996
rect 18104 6944 18110 6996
rect 21266 6944 21272 6996
rect 21324 6944 21330 6996
rect 22462 6944 22468 6996
rect 22520 6944 22526 6996
rect 25406 6944 25412 6996
rect 25464 6944 25470 6996
rect 26602 6984 26608 6996
rect 26436 6956 26608 6984
rect 11146 6876 11152 6928
rect 11204 6916 11210 6928
rect 11204 6888 12434 6916
rect 11204 6876 11210 6888
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4614 6848 4620 6860
rect 4295 6820 4620 6848
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 4614 6808 4620 6820
rect 4672 6848 4678 6860
rect 5074 6848 5080 6860
rect 4672 6820 5080 6848
rect 4672 6808 4678 6820
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 12406 6848 12434 6888
rect 17310 6876 17316 6928
rect 17368 6916 17374 6928
rect 17681 6919 17739 6925
rect 17681 6916 17693 6919
rect 17368 6888 17693 6916
rect 17368 6876 17374 6888
rect 17681 6885 17693 6888
rect 17727 6916 17739 6919
rect 17727 6888 18460 6916
rect 17727 6885 17739 6888
rect 17681 6879 17739 6885
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 12406 6820 12633 6848
rect 12621 6817 12633 6820
rect 12667 6848 12679 6851
rect 13722 6848 13728 6860
rect 12667 6820 13728 6848
rect 12667 6817 12679 6820
rect 12621 6811 12679 6817
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 15473 6851 15531 6857
rect 15473 6817 15485 6851
rect 15519 6848 15531 6851
rect 15746 6848 15752 6860
rect 15519 6820 15752 6848
rect 15519 6817 15531 6820
rect 15473 6811 15531 6817
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 18432 6848 18460 6888
rect 17920 6820 18368 6848
rect 17920 6808 17926 6820
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8260 6752 8953 6780
rect 8260 6740 8266 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9490 6780 9496 6792
rect 9171 6752 9496 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 12894 6740 12900 6792
rect 12952 6740 12958 6792
rect 15194 6740 15200 6792
rect 15252 6740 15258 6792
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 17957 6783 18015 6789
rect 17957 6749 17969 6783
rect 18003 6780 18015 6783
rect 18141 6783 18199 6789
rect 18141 6780 18153 6783
rect 18003 6752 18153 6780
rect 18003 6749 18015 6752
rect 17957 6743 18015 6749
rect 18141 6749 18153 6752
rect 18187 6780 18199 6783
rect 18230 6780 18236 6792
rect 18187 6752 18236 6780
rect 18187 6749 18199 6752
rect 18141 6743 18199 6749
rect 4522 6672 4528 6724
rect 4580 6672 4586 6724
rect 6454 6712 6460 6724
rect 5750 6684 6460 6712
rect 6454 6672 6460 6684
rect 6512 6712 6518 6724
rect 6512 6684 8524 6712
rect 6512 6672 6518 6684
rect 8496 6656 8524 6684
rect 16758 6672 16764 6724
rect 16816 6672 16822 6724
rect 17604 6712 17632 6743
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 18340 6789 18368 6820
rect 18432 6820 19012 6848
rect 18432 6789 18460 6820
rect 18984 6792 19012 6820
rect 19978 6808 19984 6860
rect 20036 6808 20042 6860
rect 20441 6851 20499 6857
rect 20441 6817 20453 6851
rect 20487 6848 20499 6851
rect 21284 6848 21312 6944
rect 20487 6820 21312 6848
rect 22480 6848 22508 6944
rect 24780 6888 24992 6916
rect 24780 6848 24808 6888
rect 22480 6820 24808 6848
rect 20487 6817 20499 6820
rect 20441 6811 20499 6817
rect 24854 6808 24860 6860
rect 24912 6808 24918 6860
rect 24964 6848 24992 6888
rect 24964 6820 25728 6848
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 18417 6783 18475 6789
rect 18417 6749 18429 6783
rect 18463 6749 18475 6783
rect 18417 6743 18475 6749
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 18598 6780 18604 6792
rect 18555 6752 18604 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 18524 6712 18552 6743
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 18966 6740 18972 6792
rect 19024 6740 19030 6792
rect 20073 6783 20131 6789
rect 20073 6749 20085 6783
rect 20119 6780 20131 6783
rect 20622 6780 20628 6792
rect 20119 6752 20628 6780
rect 20119 6749 20131 6752
rect 20073 6743 20131 6749
rect 20622 6740 20628 6752
rect 20680 6740 20686 6792
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 17604 6684 18552 6712
rect 18785 6715 18843 6721
rect 18785 6681 18797 6715
rect 18831 6712 18843 6715
rect 21192 6712 21220 6743
rect 21266 6740 21272 6792
rect 21324 6740 21330 6792
rect 21358 6740 21364 6792
rect 21416 6780 21422 6792
rect 21453 6783 21511 6789
rect 21453 6780 21465 6783
rect 21416 6752 21465 6780
rect 21416 6740 21422 6752
rect 21453 6749 21465 6752
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 24946 6740 24952 6792
rect 25004 6740 25010 6792
rect 25590 6740 25596 6792
rect 25648 6740 25654 6792
rect 25700 6789 25728 6820
rect 25792 6820 26372 6848
rect 25685 6783 25743 6789
rect 25685 6749 25697 6783
rect 25731 6749 25743 6783
rect 25685 6743 25743 6749
rect 22094 6712 22100 6724
rect 18831 6684 22100 6712
rect 18831 6681 18843 6684
rect 18785 6675 18843 6681
rect 22094 6672 22100 6684
rect 22152 6672 22158 6724
rect 25406 6672 25412 6724
rect 25464 6712 25470 6724
rect 25792 6712 25820 6820
rect 25961 6783 26019 6789
rect 25961 6749 25973 6783
rect 26007 6780 26019 6783
rect 26050 6780 26056 6792
rect 26007 6752 26056 6780
rect 26007 6749 26019 6752
rect 25961 6743 26019 6749
rect 26050 6740 26056 6752
rect 26108 6740 26114 6792
rect 26145 6783 26203 6789
rect 26145 6749 26157 6783
rect 26191 6749 26203 6783
rect 26145 6743 26203 6749
rect 25464 6684 25820 6712
rect 26160 6712 26188 6743
rect 26234 6740 26240 6792
rect 26292 6740 26298 6792
rect 26344 6789 26372 6820
rect 26329 6783 26387 6789
rect 26329 6749 26341 6783
rect 26375 6749 26387 6783
rect 26329 6743 26387 6749
rect 26436 6712 26464 6956
rect 26602 6944 26608 6956
rect 26660 6944 26666 6996
rect 28718 6944 28724 6996
rect 28776 6984 28782 6996
rect 28902 6984 28908 6996
rect 28776 6956 28908 6984
rect 28776 6944 28782 6956
rect 28902 6944 28908 6956
rect 28960 6984 28966 6996
rect 30926 6984 30932 6996
rect 28960 6956 30932 6984
rect 28960 6944 28966 6956
rect 30926 6944 30932 6956
rect 30984 6944 30990 6996
rect 31294 6944 31300 6996
rect 31352 6944 31358 6996
rect 31386 6944 31392 6996
rect 31444 6984 31450 6996
rect 31481 6987 31539 6993
rect 31481 6984 31493 6987
rect 31444 6956 31493 6984
rect 31444 6944 31450 6956
rect 31481 6953 31493 6956
rect 31527 6953 31539 6987
rect 31481 6947 31539 6953
rect 27065 6919 27123 6925
rect 27065 6916 27077 6919
rect 26620 6888 27077 6916
rect 26620 6848 26648 6888
rect 27065 6885 27077 6888
rect 27111 6885 27123 6919
rect 27065 6879 27123 6885
rect 27890 6876 27896 6928
rect 27948 6916 27954 6928
rect 30653 6919 30711 6925
rect 27948 6888 28994 6916
rect 27948 6876 27954 6888
rect 28460 6860 28488 6888
rect 26160 6684 26464 6712
rect 26528 6820 26648 6848
rect 27249 6851 27307 6857
rect 25464 6672 25470 6684
rect 8478 6604 8484 6656
rect 8536 6604 8542 6656
rect 9030 6604 9036 6656
rect 9088 6604 9094 6656
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14553 6647 14611 6653
rect 14553 6644 14565 6647
rect 13872 6616 14565 6644
rect 13872 6604 13878 6616
rect 14553 6613 14565 6616
rect 14599 6613 14611 6647
rect 14553 6607 14611 6613
rect 21637 6647 21695 6653
rect 21637 6613 21649 6647
rect 21683 6644 21695 6647
rect 22370 6644 22376 6656
rect 21683 6616 22376 6644
rect 21683 6613 21695 6616
rect 21637 6607 21695 6613
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 25314 6604 25320 6656
rect 25372 6604 25378 6656
rect 25590 6604 25596 6656
rect 25648 6644 25654 6656
rect 26528 6644 26556 6820
rect 27249 6817 27261 6851
rect 27295 6848 27307 6851
rect 27798 6848 27804 6860
rect 27295 6820 27804 6848
rect 27295 6817 27307 6820
rect 27249 6811 27307 6817
rect 27798 6808 27804 6820
rect 27856 6808 27862 6860
rect 27908 6820 28212 6848
rect 26970 6740 26976 6792
rect 27028 6740 27034 6792
rect 27525 6783 27583 6789
rect 27525 6749 27537 6783
rect 27571 6749 27583 6783
rect 27525 6743 27583 6749
rect 27618 6783 27676 6789
rect 27618 6749 27630 6783
rect 27664 6780 27676 6783
rect 27706 6780 27712 6792
rect 27664 6752 27712 6780
rect 27664 6749 27676 6752
rect 27618 6743 27676 6749
rect 27249 6715 27307 6721
rect 27249 6681 27261 6715
rect 27295 6712 27307 6715
rect 27547 6712 27575 6743
rect 27706 6740 27712 6752
rect 27764 6740 27770 6792
rect 27908 6789 27936 6820
rect 28184 6792 28212 6820
rect 28442 6808 28448 6860
rect 28500 6808 28506 6860
rect 28534 6808 28540 6860
rect 28592 6808 28598 6860
rect 28966 6848 28994 6888
rect 30653 6885 30665 6919
rect 30699 6916 30711 6919
rect 31312 6916 31340 6944
rect 30699 6888 31340 6916
rect 30699 6885 30711 6888
rect 30653 6879 30711 6885
rect 32493 6851 32551 6857
rect 32493 6848 32505 6851
rect 28966 6820 32505 6848
rect 32493 6817 32505 6820
rect 32539 6817 32551 6851
rect 32493 6811 32551 6817
rect 32582 6808 32588 6860
rect 32640 6808 32646 6860
rect 32858 6808 32864 6860
rect 32916 6848 32922 6860
rect 32953 6851 33011 6857
rect 32953 6848 32965 6851
rect 32916 6820 32965 6848
rect 32916 6808 32922 6820
rect 32953 6817 32965 6820
rect 32999 6817 33011 6851
rect 32953 6811 33011 6817
rect 33134 6808 33140 6860
rect 33192 6808 33198 6860
rect 27893 6783 27951 6789
rect 27893 6749 27905 6783
rect 27939 6749 27951 6783
rect 27893 6743 27951 6749
rect 27982 6740 27988 6792
rect 28040 6789 28046 6792
rect 28040 6743 28048 6789
rect 28040 6740 28046 6743
rect 28166 6740 28172 6792
rect 28224 6740 28230 6792
rect 28258 6740 28264 6792
rect 28316 6740 28322 6792
rect 28353 6783 28411 6789
rect 28353 6749 28365 6783
rect 28399 6749 28411 6783
rect 28353 6743 28411 6749
rect 27295 6684 27575 6712
rect 27801 6715 27859 6721
rect 27295 6681 27307 6684
rect 27249 6675 27307 6681
rect 27801 6681 27813 6715
rect 27847 6712 27859 6715
rect 28074 6712 28080 6724
rect 27847 6684 28080 6712
rect 27847 6681 27859 6684
rect 27801 6675 27859 6681
rect 28074 6672 28080 6684
rect 28132 6672 28138 6724
rect 28368 6712 28396 6743
rect 28718 6740 28724 6792
rect 28776 6740 28782 6792
rect 28810 6740 28816 6792
rect 28868 6780 28874 6792
rect 29917 6783 29975 6789
rect 29917 6780 29929 6783
rect 28868 6752 29929 6780
rect 28868 6740 28874 6752
rect 29917 6749 29929 6752
rect 29963 6749 29975 6783
rect 29917 6743 29975 6749
rect 30101 6783 30159 6789
rect 30101 6749 30113 6783
rect 30147 6749 30159 6783
rect 30101 6743 30159 6749
rect 30377 6783 30435 6789
rect 30377 6749 30389 6783
rect 30423 6780 30435 6783
rect 30466 6780 30472 6792
rect 30423 6752 30472 6780
rect 30423 6749 30435 6752
rect 30377 6743 30435 6749
rect 28184 6684 28396 6712
rect 25648 6616 26556 6644
rect 26605 6647 26663 6653
rect 25648 6604 25654 6616
rect 26605 6613 26617 6647
rect 26651 6644 26663 6647
rect 27430 6644 27436 6656
rect 26651 6616 27436 6644
rect 26651 6613 26663 6616
rect 26605 6607 26663 6613
rect 27430 6604 27436 6616
rect 27488 6604 27494 6656
rect 28184 6653 28212 6684
rect 28169 6647 28227 6653
rect 28169 6613 28181 6647
rect 28215 6613 28227 6647
rect 28169 6607 28227 6613
rect 28350 6604 28356 6656
rect 28408 6644 28414 6656
rect 30116 6644 30144 6743
rect 30466 6740 30472 6752
rect 30524 6740 30530 6792
rect 30558 6740 30564 6792
rect 30616 6780 30622 6792
rect 30745 6783 30803 6789
rect 30745 6780 30757 6783
rect 30616 6752 30757 6780
rect 30616 6740 30622 6752
rect 30745 6749 30757 6752
rect 30791 6749 30803 6783
rect 30745 6743 30803 6749
rect 30834 6740 30840 6792
rect 30892 6740 30898 6792
rect 31754 6740 31760 6792
rect 31812 6740 31818 6792
rect 31849 6783 31907 6789
rect 31849 6749 31861 6783
rect 31895 6749 31907 6783
rect 31849 6743 31907 6749
rect 31941 6783 31999 6789
rect 31941 6749 31953 6783
rect 31987 6749 31999 6783
rect 31941 6743 31999 6749
rect 28408 6616 30144 6644
rect 31864 6644 31892 6743
rect 31956 6712 31984 6743
rect 32122 6740 32128 6792
rect 32180 6740 32186 6792
rect 32674 6740 32680 6792
rect 32732 6740 32738 6792
rect 32769 6783 32827 6789
rect 32769 6749 32781 6783
rect 32815 6749 32827 6783
rect 32769 6743 32827 6749
rect 32784 6712 32812 6743
rect 33042 6740 33048 6792
rect 33100 6780 33106 6792
rect 33229 6783 33287 6789
rect 33229 6780 33241 6783
rect 33100 6752 33241 6780
rect 33100 6740 33106 6752
rect 33229 6749 33241 6752
rect 33275 6749 33287 6783
rect 33229 6743 33287 6749
rect 31956 6684 32812 6712
rect 32232 6656 32260 6684
rect 34422 6672 34428 6724
rect 34480 6672 34486 6724
rect 31938 6644 31944 6656
rect 31864 6616 31944 6644
rect 28408 6604 28414 6616
rect 31938 6604 31944 6616
rect 31996 6604 32002 6656
rect 32214 6604 32220 6656
rect 32272 6604 32278 6656
rect 33597 6647 33655 6653
rect 33597 6613 33609 6647
rect 33643 6644 33655 6647
rect 34440 6644 34468 6672
rect 33643 6616 34468 6644
rect 33643 6613 33655 6616
rect 33597 6607 33655 6613
rect 1104 6554 38272 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38272 6554
rect 1104 6480 38272 6502
rect 4522 6400 4528 6452
rect 4580 6440 4586 6452
rect 4709 6443 4767 6449
rect 4709 6440 4721 6443
rect 4580 6412 4721 6440
rect 4580 6400 4586 6412
rect 4709 6409 4721 6412
rect 4755 6409 4767 6443
rect 4709 6403 4767 6409
rect 5166 6400 5172 6452
rect 5224 6400 5230 6452
rect 7837 6443 7895 6449
rect 7837 6409 7849 6443
rect 7883 6440 7895 6443
rect 9490 6440 9496 6452
rect 7883 6412 9496 6440
rect 7883 6409 7895 6412
rect 7837 6403 7895 6409
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 13906 6400 13912 6452
rect 13964 6440 13970 6452
rect 14277 6443 14335 6449
rect 14277 6440 14289 6443
rect 13964 6412 14289 6440
rect 13964 6400 13970 6412
rect 14277 6409 14289 6412
rect 14323 6409 14335 6443
rect 14277 6403 14335 6409
rect 15289 6443 15347 6449
rect 15289 6409 15301 6443
rect 15335 6409 15347 6443
rect 15289 6403 15347 6409
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6304 4951 6307
rect 5184 6304 5212 6400
rect 7745 6375 7803 6381
rect 7745 6341 7757 6375
rect 7791 6372 7803 6375
rect 8846 6372 8852 6384
rect 7791 6344 8852 6372
rect 7791 6341 7803 6344
rect 7745 6335 7803 6341
rect 8846 6332 8852 6344
rect 8904 6332 8910 6384
rect 9398 6332 9404 6384
rect 9456 6372 9462 6384
rect 9953 6375 10011 6381
rect 9953 6372 9965 6375
rect 9456 6344 9965 6372
rect 9456 6332 9462 6344
rect 9953 6341 9965 6344
rect 9999 6341 10011 6375
rect 14642 6372 14648 6384
rect 9953 6335 10011 6341
rect 14568 6344 14648 6372
rect 4939 6276 5212 6304
rect 4939 6273 4951 6276
rect 4893 6267 4951 6273
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8389 6307 8447 6313
rect 8389 6304 8401 6307
rect 8260 6276 8401 6304
rect 8260 6264 8266 6276
rect 8389 6273 8401 6276
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6304 9735 6307
rect 10045 6307 10103 6313
rect 10045 6304 10057 6307
rect 9723 6276 10057 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 10045 6273 10057 6276
rect 10091 6304 10103 6307
rect 10226 6304 10232 6316
rect 10091 6276 10232 6304
rect 10091 6273 10103 6276
rect 10045 6267 10103 6273
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 7524 6208 7941 6236
rect 7524 6196 7530 6208
rect 7929 6205 7941 6208
rect 7975 6236 7987 6239
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 7975 6208 8585 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8573 6205 8585 6208
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6236 8723 6239
rect 8757 6239 8815 6245
rect 8757 6236 8769 6239
rect 8711 6208 8769 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 8757 6205 8769 6208
rect 8803 6205 8815 6239
rect 8757 6199 8815 6205
rect 8588 6168 8616 6199
rect 9306 6196 9312 6248
rect 9364 6196 9370 6248
rect 9508 6236 9536 6267
rect 10226 6264 10232 6276
rect 10284 6304 10290 6316
rect 12253 6307 12311 6313
rect 12253 6304 12265 6307
rect 10284 6276 12265 6304
rect 10284 6264 10290 6276
rect 12253 6273 12265 6276
rect 12299 6273 12311 6307
rect 12253 6267 12311 6273
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12529 6307 12587 6313
rect 12529 6304 12541 6307
rect 12483 6276 12541 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12529 6273 12541 6276
rect 12575 6273 12587 6307
rect 12529 6267 12587 6273
rect 12805 6307 12863 6313
rect 12805 6273 12817 6307
rect 12851 6304 12863 6307
rect 13630 6304 13636 6316
rect 12851 6276 13636 6304
rect 12851 6273 12863 6276
rect 12805 6267 12863 6273
rect 9766 6236 9772 6248
rect 9508 6208 9772 6236
rect 9766 6196 9772 6208
rect 9824 6236 9830 6248
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 9824 6208 12081 6236
rect 9824 6196 9830 6208
rect 12069 6205 12081 6208
rect 12115 6205 12127 6239
rect 12268 6236 12296 6267
rect 13630 6264 13636 6276
rect 13688 6264 13694 6316
rect 14568 6313 14596 6344
rect 14642 6332 14648 6344
rect 14700 6372 14706 6384
rect 15304 6372 15332 6403
rect 17862 6400 17868 6452
rect 17920 6400 17926 6452
rect 18690 6400 18696 6452
rect 18748 6400 18754 6452
rect 19334 6400 19340 6452
rect 19392 6400 19398 6452
rect 19889 6443 19947 6449
rect 19889 6409 19901 6443
rect 19935 6440 19947 6443
rect 19978 6440 19984 6452
rect 19935 6412 19984 6440
rect 19935 6409 19947 6412
rect 19889 6403 19947 6409
rect 19978 6400 19984 6412
rect 20036 6400 20042 6452
rect 20070 6400 20076 6452
rect 20128 6400 20134 6452
rect 23290 6400 23296 6452
rect 23348 6440 23354 6452
rect 23753 6443 23811 6449
rect 23348 6412 23520 6440
rect 23348 6400 23354 6412
rect 14700 6344 15332 6372
rect 17880 6372 17908 6400
rect 17880 6344 18276 6372
rect 14700 6332 14706 6344
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 15013 6307 15071 6313
rect 15013 6273 15025 6307
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 12618 6236 12624 6248
rect 12268 6208 12624 6236
rect 12069 6199 12127 6205
rect 9677 6171 9735 6177
rect 9677 6168 9689 6171
rect 8588 6140 9689 6168
rect 9677 6137 9689 6140
rect 9723 6137 9735 6171
rect 12084 6168 12112 6199
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 12342 6168 12348 6180
rect 12084 6140 12348 6168
rect 9677 6131 9735 6137
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 7374 6060 7380 6112
rect 7432 6060 7438 6112
rect 8202 6060 8208 6112
rect 8260 6060 8266 6112
rect 8846 6060 8852 6112
rect 8904 6100 8910 6112
rect 9490 6100 9496 6112
rect 8904 6072 9496 6100
rect 8904 6060 8910 6072
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 14844 6100 14872 6199
rect 15028 6168 15056 6267
rect 15286 6264 15292 6316
rect 15344 6264 15350 6316
rect 15378 6264 15384 6316
rect 15436 6264 15442 6316
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6304 18107 6307
rect 18138 6304 18144 6316
rect 18095 6276 18144 6304
rect 18095 6273 18107 6276
rect 18049 6267 18107 6273
rect 15304 6236 15332 6264
rect 15580 6236 15608 6267
rect 18138 6264 18144 6276
rect 18196 6264 18202 6316
rect 18248 6313 18276 6344
rect 18598 6332 18604 6384
rect 18656 6372 18662 6384
rect 19061 6375 19119 6381
rect 19061 6372 19073 6375
rect 18656 6344 19073 6372
rect 18656 6332 18662 6344
rect 19061 6341 19073 6344
rect 19107 6341 19119 6375
rect 19061 6335 19119 6341
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 18325 6307 18383 6313
rect 18325 6273 18337 6307
rect 18371 6273 18383 6307
rect 18325 6267 18383 6273
rect 18509 6307 18567 6313
rect 18509 6273 18521 6307
rect 18555 6304 18567 6307
rect 18616 6304 18644 6332
rect 18555 6276 18644 6304
rect 18877 6307 18935 6313
rect 18555 6273 18567 6276
rect 18509 6267 18567 6273
rect 18877 6273 18889 6307
rect 18923 6304 18935 6307
rect 18966 6304 18972 6316
rect 18923 6276 18972 6304
rect 18923 6273 18935 6276
rect 18877 6267 18935 6273
rect 15304 6208 15608 6236
rect 18156 6236 18184 6264
rect 18340 6236 18368 6267
rect 18892 6236 18920 6267
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 19352 6304 19380 6400
rect 19702 6304 19708 6316
rect 19352 6276 19708 6304
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 19889 6307 19947 6313
rect 19889 6273 19901 6307
rect 19935 6304 19947 6307
rect 20088 6304 20116 6400
rect 22373 6375 22431 6381
rect 22373 6341 22385 6375
rect 22419 6372 22431 6375
rect 22554 6372 22560 6384
rect 22419 6344 22560 6372
rect 22419 6341 22431 6344
rect 22373 6335 22431 6341
rect 22554 6332 22560 6344
rect 22612 6332 22618 6384
rect 22922 6332 22928 6384
rect 22980 6372 22986 6384
rect 23492 6381 23520 6412
rect 23753 6409 23765 6443
rect 23799 6409 23811 6443
rect 23753 6403 23811 6409
rect 24219 6443 24277 6449
rect 24219 6409 24231 6443
rect 24265 6440 24277 6443
rect 24946 6440 24952 6452
rect 24265 6412 24952 6440
rect 24265 6409 24277 6412
rect 24219 6403 24277 6409
rect 23385 6375 23443 6381
rect 23385 6372 23397 6375
rect 22980 6344 23397 6372
rect 22980 6332 22986 6344
rect 23385 6341 23397 6344
rect 23431 6341 23443 6375
rect 23385 6335 23443 6341
rect 23477 6375 23535 6381
rect 23477 6341 23489 6375
rect 23523 6341 23535 6375
rect 23768 6372 23796 6403
rect 24946 6400 24952 6412
rect 25004 6400 25010 6452
rect 25222 6400 25228 6452
rect 25280 6440 25286 6452
rect 25501 6443 25559 6449
rect 25501 6440 25513 6443
rect 25280 6412 25513 6440
rect 25280 6400 25286 6412
rect 25501 6409 25513 6412
rect 25547 6409 25559 6443
rect 25501 6403 25559 6409
rect 27982 6400 27988 6452
rect 28040 6400 28046 6452
rect 28166 6400 28172 6452
rect 28224 6440 28230 6452
rect 31018 6440 31024 6452
rect 28224 6412 31024 6440
rect 28224 6400 28230 6412
rect 31018 6400 31024 6412
rect 31076 6400 31082 6452
rect 33134 6440 33140 6452
rect 31726 6412 33140 6440
rect 24121 6375 24179 6381
rect 24121 6372 24133 6375
rect 23768 6344 24133 6372
rect 23477 6335 23535 6341
rect 24121 6341 24133 6344
rect 24167 6341 24179 6375
rect 24121 6335 24179 6341
rect 24486 6332 24492 6384
rect 24544 6372 24550 6384
rect 24544 6344 25268 6372
rect 24544 6332 24550 6344
rect 19935 6276 20116 6304
rect 19935 6273 19947 6276
rect 19889 6267 19947 6273
rect 18156 6208 18368 6236
rect 18616 6208 18920 6236
rect 15028 6140 15424 6168
rect 15396 6112 15424 6140
rect 18138 6128 18144 6180
rect 18196 6128 18202 6180
rect 15194 6100 15200 6112
rect 14844 6072 15200 6100
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15378 6060 15384 6112
rect 15436 6060 15442 6112
rect 15657 6103 15715 6109
rect 15657 6069 15669 6103
rect 15703 6100 15715 6103
rect 16482 6100 16488 6112
rect 15703 6072 16488 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 18509 6103 18567 6109
rect 18509 6069 18521 6103
rect 18555 6100 18567 6103
rect 18616 6100 18644 6208
rect 22572 6168 22600 6332
rect 22646 6264 22652 6316
rect 22704 6264 22710 6316
rect 22741 6307 22799 6313
rect 22741 6273 22753 6307
rect 22787 6304 22799 6307
rect 23106 6304 23112 6316
rect 22787 6276 23112 6304
rect 22787 6273 22799 6276
rect 22741 6267 22799 6273
rect 23106 6264 23112 6276
rect 23164 6304 23170 6316
rect 23201 6307 23259 6313
rect 23201 6304 23213 6307
rect 23164 6276 23213 6304
rect 23164 6264 23170 6276
rect 23201 6273 23213 6276
rect 23247 6273 23259 6307
rect 23201 6267 23259 6273
rect 23566 6264 23572 6316
rect 23624 6264 23630 6316
rect 24026 6264 24032 6316
rect 24084 6304 24090 6316
rect 24305 6307 24363 6313
rect 24305 6304 24317 6307
rect 24084 6276 24317 6304
rect 24084 6264 24090 6276
rect 24305 6273 24317 6276
rect 24351 6273 24363 6307
rect 24305 6267 24363 6273
rect 24397 6307 24455 6313
rect 24397 6273 24409 6307
rect 24443 6273 24455 6307
rect 25240 6304 25268 6344
rect 25314 6332 25320 6384
rect 25372 6372 25378 6384
rect 31726 6372 31754 6412
rect 33134 6400 33140 6412
rect 33192 6400 33198 6452
rect 25372 6344 31754 6372
rect 32769 6375 32827 6381
rect 25372 6332 25378 6344
rect 32769 6341 32781 6375
rect 32815 6341 32827 6375
rect 32769 6335 32827 6341
rect 25409 6307 25467 6313
rect 25409 6304 25421 6307
rect 25240 6276 25421 6304
rect 24397 6267 24455 6273
rect 25409 6273 25421 6276
rect 25455 6273 25467 6307
rect 25409 6267 25467 6273
rect 25593 6307 25651 6313
rect 25593 6273 25605 6307
rect 25639 6304 25651 6307
rect 26050 6304 26056 6316
rect 25639 6276 26056 6304
rect 25639 6273 25651 6276
rect 25593 6267 25651 6273
rect 22664 6236 22692 6264
rect 22833 6239 22891 6245
rect 22833 6236 22845 6239
rect 22664 6208 22845 6236
rect 22833 6205 22845 6208
rect 22879 6205 22891 6239
rect 22833 6199 22891 6205
rect 24412 6180 24440 6267
rect 25424 6236 25452 6267
rect 26050 6264 26056 6276
rect 26108 6264 26114 6316
rect 27798 6304 27804 6316
rect 27356 6276 27804 6304
rect 26786 6236 26792 6248
rect 25424 6208 26792 6236
rect 26786 6196 26792 6208
rect 26844 6196 26850 6248
rect 22572 6140 23980 6168
rect 18555 6072 18644 6100
rect 19245 6103 19303 6109
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 19245 6069 19257 6103
rect 19291 6100 19303 6103
rect 19518 6100 19524 6112
rect 19291 6072 19524 6100
rect 19291 6069 19303 6072
rect 19245 6063 19303 6069
rect 19518 6060 19524 6072
rect 19576 6060 19582 6112
rect 23014 6060 23020 6112
rect 23072 6060 23078 6112
rect 23952 6100 23980 6140
rect 24394 6128 24400 6180
rect 24452 6128 24458 6180
rect 27356 6100 27384 6276
rect 27798 6264 27804 6276
rect 27856 6264 27862 6316
rect 28077 6307 28135 6313
rect 28077 6273 28089 6307
rect 28123 6273 28135 6307
rect 28077 6267 28135 6273
rect 28261 6307 28319 6313
rect 28261 6273 28273 6307
rect 28307 6273 28319 6307
rect 28261 6267 28319 6273
rect 27525 6239 27583 6245
rect 27525 6236 27537 6239
rect 27448 6208 27537 6236
rect 27448 6180 27476 6208
rect 27525 6205 27537 6208
rect 27571 6205 27583 6239
rect 27525 6199 27583 6205
rect 27614 6196 27620 6248
rect 27672 6236 27678 6248
rect 28092 6236 28120 6267
rect 27672 6208 28120 6236
rect 27672 6196 27678 6208
rect 27430 6128 27436 6180
rect 27488 6168 27494 6180
rect 28276 6168 28304 6267
rect 32214 6264 32220 6316
rect 32272 6304 32278 6316
rect 32493 6307 32551 6313
rect 32493 6304 32505 6307
rect 32272 6276 32505 6304
rect 32272 6264 32278 6276
rect 32493 6273 32505 6276
rect 32539 6273 32551 6307
rect 32493 6267 32551 6273
rect 32585 6307 32643 6313
rect 32585 6273 32597 6307
rect 32631 6304 32643 6307
rect 32674 6304 32680 6316
rect 32631 6276 32680 6304
rect 32631 6273 32643 6276
rect 32585 6267 32643 6273
rect 32600 6236 32628 6267
rect 32674 6264 32680 6276
rect 32732 6264 32738 6316
rect 32784 6236 32812 6335
rect 27488 6140 28304 6168
rect 32048 6208 32628 6236
rect 32692 6208 32812 6236
rect 27488 6128 27494 6140
rect 32048 6112 32076 6208
rect 32582 6128 32588 6180
rect 32640 6168 32646 6180
rect 32692 6168 32720 6208
rect 32640 6140 32720 6168
rect 32640 6128 32646 6140
rect 32766 6128 32772 6180
rect 32824 6128 32830 6180
rect 23952 6072 27384 6100
rect 27614 6060 27620 6112
rect 27672 6060 27678 6112
rect 27798 6060 27804 6112
rect 27856 6100 27862 6112
rect 28902 6100 28908 6112
rect 27856 6072 28908 6100
rect 27856 6060 27862 6072
rect 28902 6060 28908 6072
rect 28960 6060 28966 6112
rect 32030 6060 32036 6112
rect 32088 6060 32094 6112
rect 1104 6010 38272 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38272 6010
rect 1104 5936 38272 5958
rect 8202 5856 8208 5908
rect 8260 5856 8266 5908
rect 9306 5896 9312 5908
rect 9048 5868 9312 5896
rect 5074 5720 5080 5772
rect 5132 5760 5138 5772
rect 6914 5760 6920 5772
rect 5132 5732 6920 5760
rect 5132 5720 5138 5732
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5760 7251 5763
rect 8220 5760 8248 5856
rect 7239 5732 8248 5760
rect 8665 5763 8723 5769
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 8665 5729 8677 5763
rect 8711 5760 8723 5763
rect 9048 5760 9076 5868
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 10318 5856 10324 5908
rect 10376 5896 10382 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 10376 5868 12817 5896
rect 10376 5856 10382 5868
rect 12805 5865 12817 5868
rect 12851 5896 12863 5899
rect 14182 5896 14188 5908
rect 12851 5868 14188 5896
rect 12851 5865 12863 5868
rect 12805 5859 12863 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 15470 5856 15476 5908
rect 15528 5896 15534 5908
rect 15703 5899 15761 5905
rect 15703 5896 15715 5899
rect 15528 5868 15715 5896
rect 15528 5856 15534 5868
rect 15703 5865 15715 5868
rect 15749 5896 15761 5899
rect 16298 5896 16304 5908
rect 15749 5868 16304 5896
rect 15749 5865 15761 5868
rect 15703 5859 15761 5865
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 18138 5856 18144 5908
rect 18196 5856 18202 5908
rect 20070 5896 20076 5908
rect 19352 5868 20076 5896
rect 9125 5831 9183 5837
rect 9125 5797 9137 5831
rect 9171 5828 9183 5831
rect 9674 5828 9680 5840
rect 9171 5800 9680 5828
rect 9171 5797 9183 5800
rect 9125 5791 9183 5797
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 13538 5828 13544 5840
rect 9922 5800 13544 5828
rect 8711 5732 9076 5760
rect 8711 5729 8723 5732
rect 8665 5723 8723 5729
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 8478 5692 8484 5704
rect 8326 5664 8484 5692
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 9048 5701 9076 5732
rect 9309 5763 9367 5769
rect 9309 5729 9321 5763
rect 9355 5760 9367 5763
rect 9355 5732 9812 5760
rect 9355 5729 9367 5732
rect 9309 5723 9367 5729
rect 9784 5704 9812 5732
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 9398 5652 9404 5704
rect 9456 5652 9462 5704
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 9548 5664 9593 5692
rect 9548 5652 9554 5664
rect 9766 5652 9772 5704
rect 9824 5652 9830 5704
rect 9922 5701 9950 5800
rect 10318 5701 10324 5704
rect 9907 5695 9965 5701
rect 9907 5661 9919 5695
rect 9953 5661 9965 5695
rect 9907 5655 9965 5661
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10285 5695 10324 5701
rect 10285 5661 10297 5695
rect 10285 5655 10324 5661
rect 5353 5627 5411 5633
rect 5353 5593 5365 5627
rect 5399 5624 5411 5627
rect 5626 5624 5632 5636
rect 5399 5596 5632 5624
rect 5399 5593 5411 5596
rect 5353 5587 5411 5593
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 9677 5627 9735 5633
rect 9677 5593 9689 5627
rect 9723 5593 9735 5627
rect 10152 5624 10180 5655
rect 10318 5652 10324 5655
rect 10376 5652 10382 5704
rect 10658 5701 10686 5800
rect 13538 5788 13544 5800
rect 13596 5788 13602 5840
rect 14918 5760 14924 5772
rect 13924 5732 14924 5760
rect 10643 5695 10701 5701
rect 10643 5661 10655 5695
rect 10689 5661 10701 5695
rect 10643 5655 10701 5661
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 12529 5695 12587 5701
rect 12529 5692 12541 5695
rect 12492 5664 12541 5692
rect 12492 5652 12498 5664
rect 12529 5661 12541 5664
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 9677 5587 9735 5593
rect 9876 5596 10180 5624
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 8202 5556 8208 5568
rect 6871 5528 8208 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 9033 5559 9091 5565
rect 9033 5525 9045 5559
rect 9079 5556 9091 5559
rect 9692 5556 9720 5587
rect 9876 5568 9904 5596
rect 10410 5584 10416 5636
rect 10468 5584 10474 5636
rect 10505 5627 10563 5633
rect 10505 5593 10517 5627
rect 10551 5624 10563 5627
rect 11977 5627 12035 5633
rect 11977 5624 11989 5627
rect 10551 5596 11989 5624
rect 10551 5593 10563 5596
rect 10505 5587 10563 5593
rect 11977 5593 11989 5596
rect 12023 5593 12035 5627
rect 12544 5624 12572 5655
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 13924 5701 13952 5732
rect 14918 5720 14924 5732
rect 14976 5760 14982 5772
rect 14976 5732 15424 5760
rect 14976 5720 14982 5732
rect 12713 5695 12771 5701
rect 12713 5692 12725 5695
rect 12676 5664 12725 5692
rect 12676 5652 12682 5664
rect 12713 5661 12725 5664
rect 12759 5661 12771 5695
rect 12713 5655 12771 5661
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5661 12955 5695
rect 12897 5655 12955 5661
rect 13633 5695 13691 5701
rect 13633 5661 13645 5695
rect 13679 5661 13691 5695
rect 13633 5655 13691 5661
rect 13909 5695 13967 5701
rect 13909 5661 13921 5695
rect 13955 5661 13967 5695
rect 13909 5655 13967 5661
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5692 14795 5695
rect 15194 5692 15200 5704
rect 14783 5664 15200 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 12912 5624 12940 5655
rect 12986 5624 12992 5636
rect 12544 5596 12992 5624
rect 11977 5587 12035 5593
rect 12986 5584 12992 5596
rect 13044 5584 13050 5636
rect 13648 5624 13676 5655
rect 15194 5652 15200 5664
rect 15252 5652 15258 5704
rect 15396 5701 15424 5732
rect 15746 5720 15752 5772
rect 15804 5760 15810 5772
rect 17497 5763 17555 5769
rect 17497 5760 17509 5763
rect 15804 5732 17509 5760
rect 15804 5720 15810 5732
rect 17497 5729 17509 5732
rect 17543 5729 17555 5763
rect 17497 5723 17555 5729
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 17126 5652 17132 5704
rect 17184 5652 17190 5704
rect 18156 5692 18184 5856
rect 19352 5828 19380 5868
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 22649 5899 22707 5905
rect 22649 5865 22661 5899
rect 22695 5896 22707 5899
rect 22830 5896 22836 5908
rect 22695 5868 22836 5896
rect 22695 5865 22707 5868
rect 22649 5859 22707 5865
rect 22830 5856 22836 5868
rect 22888 5856 22894 5908
rect 23198 5856 23204 5908
rect 23256 5896 23262 5908
rect 27430 5896 27436 5908
rect 23256 5868 27436 5896
rect 23256 5856 23262 5868
rect 27430 5856 27436 5868
rect 27488 5856 27494 5908
rect 30466 5856 30472 5908
rect 30524 5856 30530 5908
rect 32030 5856 32036 5908
rect 32088 5856 32094 5908
rect 32214 5856 32220 5908
rect 32272 5856 32278 5908
rect 19260 5800 19380 5828
rect 22189 5831 22247 5837
rect 19260 5769 19288 5800
rect 22189 5797 22201 5831
rect 22235 5828 22247 5831
rect 23216 5828 23244 5856
rect 22235 5800 23244 5828
rect 22235 5797 22247 5800
rect 22189 5791 22247 5797
rect 24670 5788 24676 5840
rect 24728 5828 24734 5840
rect 28350 5828 28356 5840
rect 24728 5800 28356 5828
rect 24728 5788 24734 5800
rect 19245 5763 19303 5769
rect 19245 5729 19257 5763
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 19334 5720 19340 5772
rect 19392 5720 19398 5772
rect 19518 5720 19524 5772
rect 19576 5760 19582 5772
rect 19705 5763 19763 5769
rect 19705 5760 19717 5763
rect 19576 5732 19717 5760
rect 19576 5720 19582 5732
rect 19705 5729 19717 5732
rect 19751 5729 19763 5763
rect 24946 5760 24952 5772
rect 19705 5723 19763 5729
rect 22204 5732 22692 5760
rect 19352 5692 19380 5720
rect 19613 5695 19671 5701
rect 19613 5692 19625 5695
rect 18156 5664 19625 5692
rect 19613 5661 19625 5664
rect 19659 5661 19671 5695
rect 19613 5655 19671 5661
rect 20070 5652 20076 5704
rect 20128 5652 20134 5704
rect 20438 5652 20444 5704
rect 20496 5652 20502 5704
rect 20530 5652 20536 5704
rect 20588 5692 20594 5704
rect 22204 5701 22232 5732
rect 22664 5704 22692 5732
rect 24596 5732 24952 5760
rect 20625 5695 20683 5701
rect 20625 5692 20637 5695
rect 20588 5664 20637 5692
rect 20588 5652 20594 5664
rect 20625 5661 20637 5664
rect 20671 5661 20683 5695
rect 20625 5655 20683 5661
rect 22189 5695 22247 5701
rect 22189 5661 22201 5695
rect 22235 5661 22247 5695
rect 22189 5655 22247 5661
rect 22373 5695 22431 5701
rect 22373 5661 22385 5695
rect 22419 5661 22431 5695
rect 22373 5655 22431 5661
rect 14274 5624 14280 5636
rect 13648 5596 14280 5624
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 15473 5627 15531 5633
rect 15473 5593 15485 5627
rect 15519 5624 15531 5627
rect 15930 5624 15936 5636
rect 15519 5596 15936 5624
rect 15519 5593 15531 5596
rect 15473 5587 15531 5593
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 16114 5584 16120 5636
rect 16172 5584 16178 5636
rect 19337 5627 19395 5633
rect 19337 5593 19349 5627
rect 19383 5624 19395 5627
rect 19702 5624 19708 5636
rect 19383 5596 19708 5624
rect 19383 5593 19395 5596
rect 19337 5587 19395 5593
rect 19702 5584 19708 5596
rect 19760 5584 19766 5636
rect 22388 5624 22416 5655
rect 22646 5652 22652 5704
rect 22704 5652 22710 5704
rect 22922 5652 22928 5704
rect 22980 5652 22986 5704
rect 23106 5652 23112 5704
rect 23164 5652 23170 5704
rect 23566 5652 23572 5704
rect 23624 5652 23630 5704
rect 23658 5652 23664 5704
rect 23716 5652 23722 5704
rect 24394 5652 24400 5704
rect 24452 5652 24458 5704
rect 24596 5701 24624 5732
rect 24946 5720 24952 5732
rect 25004 5720 25010 5772
rect 25056 5701 25084 5800
rect 28350 5788 28356 5800
rect 28408 5788 28414 5840
rect 29270 5788 29276 5840
rect 29328 5828 29334 5840
rect 29825 5831 29883 5837
rect 29825 5828 29837 5831
rect 29328 5800 29837 5828
rect 29328 5788 29334 5800
rect 29825 5797 29837 5800
rect 29871 5797 29883 5831
rect 29825 5791 29883 5797
rect 29178 5720 29184 5772
rect 29236 5760 29242 5772
rect 29549 5763 29607 5769
rect 29549 5760 29561 5763
rect 29236 5732 29561 5760
rect 29236 5720 29242 5732
rect 29549 5729 29561 5732
rect 29595 5729 29607 5763
rect 29549 5723 29607 5729
rect 24581 5695 24639 5701
rect 24581 5661 24593 5695
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 25041 5695 25099 5701
rect 25041 5661 25053 5695
rect 25087 5661 25099 5695
rect 25041 5655 25099 5661
rect 23124 5624 23152 5652
rect 24412 5624 24440 5652
rect 24872 5624 24900 5655
rect 31754 5652 31760 5704
rect 31812 5692 31818 5704
rect 31849 5695 31907 5701
rect 31849 5692 31861 5695
rect 31812 5664 31861 5692
rect 31812 5652 31818 5664
rect 31849 5661 31861 5664
rect 31895 5661 31907 5695
rect 31849 5655 31907 5661
rect 32122 5652 32128 5704
rect 32180 5652 32186 5704
rect 32309 5695 32367 5701
rect 32309 5661 32321 5695
rect 32355 5661 32367 5695
rect 32309 5655 32367 5661
rect 22388 5596 23152 5624
rect 24320 5596 24900 5624
rect 30101 5627 30159 5633
rect 9079 5528 9720 5556
rect 9079 5525 9091 5528
rect 9033 5519 9091 5525
rect 9858 5516 9864 5568
rect 9916 5516 9922 5568
rect 10042 5516 10048 5568
rect 10100 5516 10106 5568
rect 10781 5559 10839 5565
rect 10781 5525 10793 5559
rect 10827 5556 10839 5559
rect 11698 5556 11704 5568
rect 10827 5528 11704 5556
rect 10827 5525 10839 5528
rect 10781 5519 10839 5525
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 13449 5559 13507 5565
rect 13449 5525 13461 5559
rect 13495 5556 13507 5559
rect 13630 5556 13636 5568
rect 13495 5528 13636 5556
rect 13495 5525 13507 5528
rect 13449 5519 13507 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 13814 5516 13820 5568
rect 13872 5516 13878 5568
rect 14366 5516 14372 5568
rect 14424 5516 14430 5568
rect 14829 5559 14887 5565
rect 14829 5525 14841 5559
rect 14875 5556 14887 5559
rect 15378 5556 15384 5568
rect 14875 5528 15384 5556
rect 14875 5525 14887 5528
rect 14829 5519 14887 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 19889 5559 19947 5565
rect 19889 5525 19901 5559
rect 19935 5556 19947 5559
rect 19978 5556 19984 5568
rect 19935 5528 19984 5556
rect 19935 5525 19947 5528
rect 19889 5519 19947 5525
rect 19978 5516 19984 5528
rect 20036 5516 20042 5568
rect 20441 5559 20499 5565
rect 20441 5525 20453 5559
rect 20487 5556 20499 5559
rect 20990 5556 20996 5568
rect 20487 5528 20996 5556
rect 20487 5525 20499 5528
rect 20441 5519 20499 5525
rect 20990 5516 20996 5528
rect 21048 5516 21054 5568
rect 22830 5516 22836 5568
rect 22888 5556 22894 5568
rect 24320 5556 24348 5596
rect 30101 5593 30113 5627
rect 30147 5624 30159 5627
rect 30190 5624 30196 5636
rect 30147 5596 30196 5624
rect 30147 5593 30159 5596
rect 30101 5587 30159 5593
rect 30190 5584 30196 5596
rect 30248 5584 30254 5636
rect 30282 5584 30288 5636
rect 30340 5584 30346 5636
rect 31665 5627 31723 5633
rect 31665 5593 31677 5627
rect 31711 5593 31723 5627
rect 31665 5587 31723 5593
rect 22888 5528 24348 5556
rect 22888 5516 22894 5528
rect 24394 5516 24400 5568
rect 24452 5516 24458 5568
rect 29822 5516 29828 5568
rect 29880 5556 29886 5568
rect 30009 5559 30067 5565
rect 30009 5556 30021 5559
rect 29880 5528 30021 5556
rect 29880 5516 29886 5528
rect 30009 5525 30021 5528
rect 30055 5556 30067 5559
rect 31680 5556 31708 5587
rect 31938 5584 31944 5636
rect 31996 5624 32002 5636
rect 32324 5624 32352 5655
rect 31996 5596 32352 5624
rect 31996 5584 32002 5596
rect 30055 5528 31708 5556
rect 30055 5525 30067 5528
rect 30009 5519 30067 5525
rect 1104 5466 38272 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38272 5466
rect 1104 5392 38272 5414
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 5684 5324 6469 5352
rect 5684 5312 5690 5324
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 7374 5312 7380 5364
rect 7432 5312 7438 5364
rect 8846 5312 8852 5364
rect 8904 5312 8910 5364
rect 9858 5352 9864 5364
rect 9324 5324 9864 5352
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 7392 5216 7420 5312
rect 6687 5188 7420 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 8202 5176 8208 5228
rect 8260 5176 8266 5228
rect 9030 5176 9036 5228
rect 9088 5216 9094 5228
rect 9324 5225 9352 5324
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 11514 5312 11520 5364
rect 11572 5352 11578 5364
rect 12158 5352 12164 5364
rect 11572 5324 12164 5352
rect 11572 5312 11578 5324
rect 12158 5312 12164 5324
rect 12216 5352 12222 5364
rect 12216 5324 13492 5352
rect 12216 5312 12222 5324
rect 9493 5287 9551 5293
rect 9493 5253 9505 5287
rect 9539 5284 9551 5287
rect 9677 5287 9735 5293
rect 9677 5284 9689 5287
rect 9539 5256 9689 5284
rect 9539 5253 9551 5256
rect 9493 5247 9551 5253
rect 9677 5253 9689 5256
rect 9723 5253 9735 5287
rect 10410 5284 10416 5296
rect 9677 5247 9735 5253
rect 9968 5256 10416 5284
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 9088 5188 9321 5216
rect 9088 5176 9094 5188
rect 9309 5185 9321 5188
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 9585 5219 9643 5225
rect 9585 5185 9597 5219
rect 9631 5216 9643 5219
rect 9858 5216 9864 5228
rect 9631 5188 9864 5216
rect 9631 5185 9643 5188
rect 9585 5179 9643 5185
rect 9858 5176 9864 5188
rect 9916 5216 9922 5228
rect 9968 5216 9996 5256
rect 10410 5244 10416 5256
rect 10468 5244 10474 5296
rect 9916 5188 9996 5216
rect 9916 5176 9922 5188
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 11532 5225 11560 5312
rect 11698 5244 11704 5296
rect 11756 5284 11762 5296
rect 11793 5287 11851 5293
rect 11793 5284 11805 5287
rect 11756 5256 11805 5284
rect 11756 5244 11762 5256
rect 11793 5253 11805 5256
rect 11839 5253 11851 5287
rect 11793 5247 11851 5253
rect 12526 5244 12532 5296
rect 12584 5244 12590 5296
rect 13464 5225 13492 5324
rect 15194 5312 15200 5364
rect 15252 5312 15258 5364
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17313 5355 17371 5361
rect 17313 5352 17325 5355
rect 17184 5324 17325 5352
rect 17184 5312 17190 5324
rect 17313 5321 17325 5324
rect 17359 5321 17371 5355
rect 17313 5315 17371 5321
rect 19705 5355 19763 5361
rect 19705 5321 19717 5355
rect 19751 5352 19763 5355
rect 20162 5352 20168 5364
rect 19751 5324 20168 5352
rect 19751 5321 19763 5324
rect 19705 5315 19763 5321
rect 20162 5312 20168 5324
rect 20220 5352 20226 5364
rect 20438 5352 20444 5364
rect 20220 5324 20444 5352
rect 20220 5312 20226 5324
rect 20438 5312 20444 5324
rect 20496 5312 20502 5364
rect 21269 5355 21327 5361
rect 21269 5321 21281 5355
rect 21315 5352 21327 5355
rect 22830 5352 22836 5364
rect 21315 5324 22836 5352
rect 21315 5321 21327 5324
rect 21269 5315 21327 5321
rect 22830 5312 22836 5324
rect 22888 5312 22894 5364
rect 23109 5355 23167 5361
rect 23109 5321 23121 5355
rect 23155 5352 23167 5355
rect 23566 5352 23572 5364
rect 23155 5324 23572 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23566 5312 23572 5324
rect 23624 5312 23630 5364
rect 23658 5312 23664 5364
rect 23716 5312 23722 5364
rect 24854 5312 24860 5364
rect 24912 5352 24918 5364
rect 27525 5355 27583 5361
rect 24912 5324 27476 5352
rect 24912 5312 24918 5324
rect 13630 5244 13636 5296
rect 13688 5284 13694 5296
rect 13725 5287 13783 5293
rect 13725 5284 13737 5287
rect 13688 5256 13737 5284
rect 13688 5244 13694 5256
rect 13725 5253 13737 5256
rect 13771 5253 13783 5287
rect 13725 5247 13783 5253
rect 19334 5244 19340 5296
rect 19392 5244 19398 5296
rect 19426 5244 19432 5296
rect 19484 5284 19490 5296
rect 19521 5287 19579 5293
rect 19521 5284 19533 5287
rect 19484 5256 19533 5284
rect 19484 5244 19490 5256
rect 19521 5253 19533 5256
rect 19567 5284 19579 5287
rect 19567 5256 20024 5284
rect 19567 5253 19579 5256
rect 19521 5247 19579 5253
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 10100 5188 10517 5216
rect 10100 5176 10106 5188
rect 10505 5185 10517 5188
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 13449 5219 13507 5225
rect 13449 5185 13461 5219
rect 13495 5185 13507 5219
rect 16114 5216 16120 5228
rect 13449 5179 13507 5185
rect 14752 5188 16120 5216
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10229 5151 10287 5157
rect 10229 5148 10241 5151
rect 9732 5120 10241 5148
rect 9732 5108 9738 5120
rect 10229 5117 10241 5120
rect 10275 5117 10287 5151
rect 10229 5111 10287 5117
rect 12986 5108 12992 5160
rect 13044 5108 13050 5160
rect 13004 5080 13032 5108
rect 13265 5083 13323 5089
rect 13265 5080 13277 5083
rect 13004 5052 13277 5080
rect 13265 5049 13277 5052
rect 13311 5049 13323 5083
rect 13265 5043 13323 5049
rect 9122 4972 9128 5024
rect 9180 4972 9186 5024
rect 11146 4972 11152 5024
rect 11204 4972 11210 5024
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 14752 5012 14780 5188
rect 16114 5176 16120 5188
rect 16172 5176 16178 5228
rect 19352 5216 19380 5244
rect 19996 5225 20024 5256
rect 20990 5244 20996 5296
rect 21048 5284 21054 5296
rect 21085 5287 21143 5293
rect 21085 5284 21097 5287
rect 21048 5256 21097 5284
rect 21048 5244 21054 5256
rect 21085 5253 21097 5256
rect 21131 5253 21143 5287
rect 21085 5247 21143 5253
rect 22925 5287 22983 5293
rect 22925 5253 22937 5287
rect 22971 5284 22983 5287
rect 25869 5287 25927 5293
rect 22971 5256 23152 5284
rect 22971 5253 22983 5256
rect 22925 5247 22983 5253
rect 23124 5228 23152 5256
rect 23308 5256 25728 5284
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 19352 5188 19809 5216
rect 19797 5185 19809 5188
rect 19843 5185 19855 5219
rect 19797 5179 19855 5185
rect 19981 5219 20039 5225
rect 19981 5185 19993 5219
rect 20027 5185 20039 5219
rect 19981 5179 20039 5185
rect 20898 5176 20904 5228
rect 20956 5176 20962 5228
rect 22281 5219 22339 5225
rect 22281 5185 22293 5219
rect 22327 5216 22339 5219
rect 22738 5216 22744 5228
rect 22327 5188 22744 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 22738 5176 22744 5188
rect 22796 5176 22802 5228
rect 23014 5176 23020 5228
rect 23072 5176 23078 5228
rect 23106 5176 23112 5228
rect 23164 5176 23170 5228
rect 23198 5176 23204 5228
rect 23256 5176 23262 5228
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 15838 5148 15844 5160
rect 15436 5120 15844 5148
rect 15436 5108 15442 5120
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 16666 5108 16672 5160
rect 16724 5108 16730 5160
rect 22370 5108 22376 5160
rect 22428 5148 22434 5160
rect 23308 5148 23336 5256
rect 23385 5219 23443 5225
rect 23385 5185 23397 5219
rect 23431 5185 23443 5219
rect 23385 5179 23443 5185
rect 22428 5120 23336 5148
rect 22428 5108 22434 5120
rect 19889 5083 19947 5089
rect 19889 5049 19901 5083
rect 19935 5080 19947 5083
rect 23290 5080 23296 5092
rect 19935 5052 23296 5080
rect 19935 5049 19947 5052
rect 19889 5043 19947 5049
rect 23290 5040 23296 5052
rect 23348 5040 23354 5092
rect 23400 5024 23428 5179
rect 24670 5176 24676 5228
rect 24728 5216 24734 5228
rect 25406 5216 25412 5228
rect 24728 5188 25412 5216
rect 24728 5176 24734 5188
rect 25406 5176 25412 5188
rect 25464 5216 25470 5228
rect 25700 5225 25728 5256
rect 25869 5253 25881 5287
rect 25915 5284 25927 5287
rect 27448 5284 27476 5324
rect 27525 5321 27537 5355
rect 27571 5352 27583 5355
rect 27614 5352 27620 5364
rect 27571 5324 27620 5352
rect 27571 5321 27583 5324
rect 27525 5315 27583 5321
rect 27614 5312 27620 5324
rect 27672 5312 27678 5364
rect 29457 5355 29515 5361
rect 29457 5352 29469 5355
rect 28736 5324 29469 5352
rect 27893 5287 27951 5293
rect 27893 5284 27905 5287
rect 25915 5256 27200 5284
rect 27448 5256 27905 5284
rect 25915 5253 25927 5256
rect 25869 5247 25927 5253
rect 25593 5219 25651 5225
rect 25593 5216 25605 5219
rect 25464 5188 25605 5216
rect 25464 5176 25470 5188
rect 25593 5185 25605 5188
rect 25639 5185 25651 5219
rect 25593 5179 25651 5185
rect 25685 5219 25743 5225
rect 25685 5185 25697 5219
rect 25731 5216 25743 5219
rect 26234 5216 26240 5228
rect 25731 5188 26240 5216
rect 25731 5185 25743 5188
rect 25685 5179 25743 5185
rect 26234 5176 26240 5188
rect 26292 5176 26298 5228
rect 27172 5225 27200 5256
rect 27893 5253 27905 5256
rect 27939 5284 27951 5287
rect 28442 5284 28448 5296
rect 27939 5256 28448 5284
rect 27939 5253 27951 5256
rect 27893 5247 27951 5253
rect 28442 5244 28448 5256
rect 28500 5244 28506 5296
rect 27157 5219 27215 5225
rect 27157 5185 27169 5219
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27614 5176 27620 5228
rect 27672 5176 27678 5228
rect 27706 5176 27712 5228
rect 27764 5176 27770 5228
rect 28736 5225 28764 5324
rect 29457 5321 29469 5324
rect 29503 5352 29515 5355
rect 30193 5355 30251 5361
rect 29503 5324 29960 5352
rect 29503 5321 29515 5324
rect 29457 5315 29515 5321
rect 28920 5256 29868 5284
rect 28920 5225 28948 5256
rect 29840 5228 29868 5256
rect 28537 5219 28595 5225
rect 28537 5216 28549 5219
rect 28000 5188 28549 5216
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5148 23719 5151
rect 24394 5148 24400 5160
rect 23707 5120 24400 5148
rect 23707 5117 23719 5120
rect 23661 5111 23719 5117
rect 24394 5108 24400 5120
rect 24452 5108 24458 5160
rect 25869 5151 25927 5157
rect 25869 5117 25881 5151
rect 25915 5148 25927 5151
rect 25915 5120 26096 5148
rect 25915 5117 25927 5120
rect 25869 5111 25927 5117
rect 26068 5092 26096 5120
rect 26970 5108 26976 5160
rect 27028 5148 27034 5160
rect 27065 5151 27123 5157
rect 27065 5148 27077 5151
rect 27028 5120 27077 5148
rect 27028 5108 27034 5120
rect 27065 5117 27077 5120
rect 27111 5148 27123 5151
rect 28000 5148 28028 5188
rect 28537 5185 28549 5188
rect 28583 5185 28595 5219
rect 28537 5179 28595 5185
rect 28721 5219 28779 5225
rect 28721 5185 28733 5219
rect 28767 5185 28779 5219
rect 28721 5179 28779 5185
rect 28905 5219 28963 5225
rect 28905 5185 28917 5219
rect 28951 5185 28963 5219
rect 28905 5179 28963 5185
rect 28997 5219 29055 5225
rect 28997 5185 29009 5219
rect 29043 5216 29055 5219
rect 29270 5216 29276 5228
rect 29043 5188 29276 5216
rect 29043 5185 29055 5188
rect 28997 5179 29055 5185
rect 29270 5176 29276 5188
rect 29328 5176 29334 5228
rect 29549 5219 29607 5225
rect 29549 5185 29561 5219
rect 29595 5216 29607 5219
rect 29733 5219 29791 5225
rect 29595 5188 29684 5216
rect 29595 5185 29607 5188
rect 29549 5179 29607 5185
rect 27111 5120 28028 5148
rect 27111 5117 27123 5120
rect 27065 5111 27123 5117
rect 28258 5108 28264 5160
rect 28316 5108 28322 5160
rect 26050 5040 26056 5092
rect 26108 5040 26114 5092
rect 27893 5083 27951 5089
rect 27893 5049 27905 5083
rect 27939 5080 27951 5083
rect 28276 5080 28304 5108
rect 27939 5052 28304 5080
rect 27939 5049 27951 5052
rect 27893 5043 27951 5049
rect 29178 5040 29184 5092
rect 29236 5080 29242 5092
rect 29273 5083 29331 5089
rect 29273 5080 29285 5083
rect 29236 5052 29285 5080
rect 29236 5040 29242 5052
rect 29273 5049 29285 5052
rect 29319 5049 29331 5083
rect 29273 5043 29331 5049
rect 29656 5024 29684 5188
rect 29733 5185 29745 5219
rect 29779 5185 29791 5219
rect 29733 5179 29791 5185
rect 12584 4984 14780 5012
rect 12584 4972 12590 4984
rect 16390 4972 16396 5024
rect 16448 4972 16454 5024
rect 23382 4972 23388 5024
rect 23440 4972 23446 5024
rect 23477 5015 23535 5021
rect 23477 4981 23489 5015
rect 23523 5012 23535 5015
rect 24394 5012 24400 5024
rect 23523 4984 24400 5012
rect 23523 4981 23535 4984
rect 23477 4975 23535 4981
rect 24394 4972 24400 4984
rect 24452 4972 24458 5024
rect 29638 4972 29644 5024
rect 29696 4972 29702 5024
rect 29748 5012 29776 5179
rect 29822 5176 29828 5228
rect 29880 5176 29886 5228
rect 29932 5225 29960 5324
rect 30193 5321 30205 5355
rect 30239 5352 30251 5355
rect 30282 5352 30288 5364
rect 30239 5324 30288 5352
rect 30239 5321 30251 5324
rect 30193 5315 30251 5321
rect 30282 5312 30288 5324
rect 30340 5312 30346 5364
rect 31481 5355 31539 5361
rect 31481 5321 31493 5355
rect 31527 5352 31539 5355
rect 32122 5352 32128 5364
rect 31527 5324 32128 5352
rect 31527 5321 31539 5324
rect 31481 5315 31539 5321
rect 32122 5312 32128 5324
rect 32180 5312 32186 5364
rect 29917 5219 29975 5225
rect 29917 5185 29929 5219
rect 29963 5185 29975 5219
rect 29917 5179 29975 5185
rect 30009 5219 30067 5225
rect 30009 5185 30021 5219
rect 30055 5216 30067 5219
rect 30098 5216 30104 5228
rect 30055 5188 30104 5216
rect 30055 5185 30067 5188
rect 30009 5179 30067 5185
rect 29932 5148 29960 5179
rect 30098 5176 30104 5188
rect 30156 5216 30162 5228
rect 30469 5219 30527 5225
rect 30469 5216 30481 5219
rect 30156 5188 30481 5216
rect 30156 5176 30162 5188
rect 30469 5185 30481 5188
rect 30515 5185 30527 5219
rect 30469 5179 30527 5185
rect 30745 5219 30803 5225
rect 30745 5185 30757 5219
rect 30791 5216 30803 5219
rect 31113 5219 31171 5225
rect 30791 5188 31064 5216
rect 30791 5185 30803 5188
rect 30745 5179 30803 5185
rect 30561 5151 30619 5157
rect 30561 5148 30573 5151
rect 29932 5120 30573 5148
rect 30561 5117 30573 5120
rect 30607 5117 30619 5151
rect 30561 5111 30619 5117
rect 29822 5040 29828 5092
rect 29880 5040 29886 5092
rect 29932 5052 30420 5080
rect 29932 5012 29960 5052
rect 30006 5012 30012 5024
rect 29748 4984 30012 5012
rect 30006 4972 30012 4984
rect 30064 4972 30070 5024
rect 30282 4972 30288 5024
rect 30340 4972 30346 5024
rect 30392 5012 30420 5052
rect 30650 5040 30656 5092
rect 30708 5040 30714 5092
rect 30760 5012 30788 5179
rect 31036 5157 31064 5188
rect 31113 5185 31125 5219
rect 31159 5216 31171 5219
rect 31754 5216 31760 5228
rect 31159 5188 31760 5216
rect 31159 5185 31171 5188
rect 31113 5179 31171 5185
rect 31754 5176 31760 5188
rect 31812 5176 31818 5228
rect 31021 5151 31079 5157
rect 31021 5117 31033 5151
rect 31067 5117 31079 5151
rect 31021 5111 31079 5117
rect 30392 4984 30788 5012
rect 1104 4922 38272 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38272 4922
rect 1104 4848 38272 4870
rect 9858 4768 9864 4820
rect 9916 4768 9922 4820
rect 10952 4811 11010 4817
rect 10952 4777 10964 4811
rect 10998 4808 11010 4811
rect 11146 4808 11152 4820
rect 10998 4780 11152 4808
rect 10998 4777 11010 4780
rect 10952 4771 11010 4777
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 12437 4811 12495 4817
rect 12437 4777 12449 4811
rect 12483 4808 12495 4811
rect 12618 4808 12624 4820
rect 12483 4780 12624 4808
rect 12483 4777 12495 4780
rect 12437 4771 12495 4777
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 15838 4768 15844 4820
rect 15896 4808 15902 4820
rect 15933 4811 15991 4817
rect 15933 4808 15945 4811
rect 15896 4780 15945 4808
rect 15896 4768 15902 4780
rect 15933 4777 15945 4780
rect 15979 4777 15991 4811
rect 15933 4771 15991 4777
rect 16390 4768 16396 4820
rect 16448 4768 16454 4820
rect 16577 4811 16635 4817
rect 16577 4777 16589 4811
rect 16623 4808 16635 4811
rect 16666 4808 16672 4820
rect 16623 4780 16672 4808
rect 16623 4777 16635 4780
rect 16577 4771 16635 4777
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 19978 4768 19984 4820
rect 20036 4768 20042 4820
rect 20162 4768 20168 4820
rect 20220 4768 20226 4820
rect 20349 4811 20407 4817
rect 20349 4777 20361 4811
rect 20395 4808 20407 4811
rect 20898 4808 20904 4820
rect 20395 4780 20904 4808
rect 20395 4777 20407 4780
rect 20349 4771 20407 4777
rect 20898 4768 20904 4780
rect 20956 4768 20962 4820
rect 20990 4768 20996 4820
rect 21048 4808 21054 4820
rect 21048 4780 23336 4808
rect 21048 4768 21054 4780
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4672 10747 4675
rect 12158 4672 12164 4684
rect 10735 4644 12164 4672
rect 10735 4641 10747 4644
rect 10689 4635 10747 4641
rect 12158 4632 12164 4644
rect 12216 4672 12222 4684
rect 14185 4675 14243 4681
rect 14185 4672 14197 4675
rect 12216 4644 14197 4672
rect 12216 4632 12222 4644
rect 14185 4641 14197 4644
rect 14231 4641 14243 4675
rect 16408 4672 16436 4768
rect 19996 4740 20024 4768
rect 23308 4740 23336 4780
rect 23382 4768 23388 4820
rect 23440 4808 23446 4820
rect 23477 4811 23535 4817
rect 23477 4808 23489 4811
rect 23440 4780 23489 4808
rect 23440 4768 23446 4780
rect 23477 4777 23489 4780
rect 23523 4777 23535 4811
rect 23477 4771 23535 4777
rect 24394 4768 24400 4820
rect 24452 4768 24458 4820
rect 25498 4768 25504 4820
rect 25556 4808 25562 4820
rect 25685 4811 25743 4817
rect 25685 4808 25697 4811
rect 25556 4780 25697 4808
rect 25556 4768 25562 4780
rect 25685 4777 25697 4780
rect 25731 4777 25743 4811
rect 25685 4771 25743 4777
rect 26050 4768 26056 4820
rect 26108 4768 26114 4820
rect 27525 4811 27583 4817
rect 27525 4777 27537 4811
rect 27571 4808 27583 4811
rect 27614 4808 27620 4820
rect 27571 4780 27620 4808
rect 27571 4777 27583 4780
rect 27525 4771 27583 4777
rect 27614 4768 27620 4780
rect 27672 4768 27678 4820
rect 29178 4768 29184 4820
rect 29236 4808 29242 4820
rect 29641 4811 29699 4817
rect 29641 4808 29653 4811
rect 29236 4780 29653 4808
rect 29236 4768 29242 4780
rect 29641 4777 29653 4780
rect 29687 4777 29699 4811
rect 29641 4771 29699 4777
rect 30006 4768 30012 4820
rect 30064 4768 30070 4820
rect 30190 4768 30196 4820
rect 30248 4808 30254 4820
rect 30285 4811 30343 4817
rect 30285 4808 30297 4811
rect 30248 4780 30297 4808
rect 30248 4768 30254 4780
rect 30285 4777 30297 4780
rect 30331 4777 30343 4811
rect 30285 4771 30343 4777
rect 27890 4740 27896 4752
rect 19996 4712 23244 4740
rect 23308 4712 27896 4740
rect 14185 4635 14243 4641
rect 16040 4644 16436 4672
rect 19521 4675 19579 4681
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 3878 4604 3884 4616
rect 1811 4576 3884 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 3878 4564 3884 4576
rect 3936 4564 3942 4616
rect 9766 4564 9772 4616
rect 9824 4604 9830 4616
rect 10045 4607 10103 4613
rect 10045 4604 10057 4607
rect 9824 4576 10057 4604
rect 9824 4564 9830 4576
rect 10045 4573 10057 4576
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 10226 4564 10232 4616
rect 10284 4564 10290 4616
rect 15930 4564 15936 4616
rect 15988 4564 15994 4616
rect 16040 4613 16068 4644
rect 19521 4641 19533 4675
rect 19567 4672 19579 4675
rect 20254 4672 20260 4684
rect 19567 4644 20260 4672
rect 19567 4641 19579 4644
rect 19521 4635 19579 4641
rect 20254 4632 20260 4644
rect 20312 4672 20318 4684
rect 23216 4672 23244 4712
rect 27890 4700 27896 4712
rect 27948 4740 27954 4752
rect 29822 4740 29828 4752
rect 27948 4712 29828 4740
rect 27948 4700 27954 4712
rect 29822 4700 29828 4712
rect 29880 4740 29886 4752
rect 30650 4740 30656 4752
rect 29880 4712 30656 4740
rect 29880 4700 29886 4712
rect 30650 4700 30656 4712
rect 30708 4700 30714 4752
rect 20312 4644 21496 4672
rect 20312 4632 20318 4644
rect 16025 4607 16083 4613
rect 16025 4573 16037 4607
rect 16071 4573 16083 4607
rect 16025 4567 16083 4573
rect 16298 4564 16304 4616
rect 16356 4564 16362 4616
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4604 16451 4607
rect 16482 4604 16488 4616
rect 16439 4576 16488 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 20346 4604 20352 4616
rect 19475 4576 20352 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 20346 4564 20352 4576
rect 20404 4604 20410 4616
rect 21269 4607 21327 4613
rect 21269 4604 21281 4607
rect 20404 4576 21281 4604
rect 20404 4564 20410 4576
rect 21269 4573 21281 4576
rect 21315 4573 21327 4607
rect 21468 4604 21496 4644
rect 23216 4644 23433 4672
rect 21818 4604 21824 4616
rect 21468 4576 21824 4604
rect 21269 4567 21327 4573
rect 21818 4564 21824 4576
rect 21876 4564 21882 4616
rect 23216 4613 23244 4644
rect 23201 4607 23259 4613
rect 23201 4573 23213 4607
rect 23247 4573 23259 4607
rect 23405 4604 23433 4644
rect 23474 4632 23480 4684
rect 23532 4672 23538 4684
rect 24673 4675 24731 4681
rect 24673 4672 24685 4675
rect 23532 4644 24685 4672
rect 23532 4632 23538 4644
rect 24673 4641 24685 4644
rect 24719 4672 24731 4675
rect 25406 4672 25412 4684
rect 24719 4644 25176 4672
rect 24719 4641 24731 4644
rect 24673 4635 24731 4641
rect 24581 4607 24639 4613
rect 24581 4604 24593 4607
rect 23405 4576 24593 4604
rect 23201 4567 23259 4573
rect 24581 4573 24593 4576
rect 24627 4573 24639 4607
rect 24765 4607 24823 4613
rect 24765 4606 24777 4607
rect 24581 4567 24639 4573
rect 24688 4578 24777 4606
rect 934 4496 940 4548
rect 992 4536 998 4548
rect 1397 4539 1455 4545
rect 1397 4536 1409 4539
rect 992 4508 1409 4536
rect 992 4496 998 4508
rect 1397 4505 1409 4508
rect 1443 4505 1455 4539
rect 12526 4536 12532 4548
rect 12190 4508 12532 4536
rect 1397 4499 1455 4505
rect 12526 4496 12532 4508
rect 12584 4496 12590 4548
rect 14458 4496 14464 4548
rect 14516 4496 14522 4548
rect 15948 4536 15976 4564
rect 22744 4548 22796 4554
rect 16209 4539 16267 4545
rect 16209 4536 16221 4539
rect 15686 4508 15884 4536
rect 15948 4508 16221 4536
rect 15856 4468 15884 4508
rect 16209 4505 16221 4508
rect 16255 4505 16267 4539
rect 19981 4539 20039 4545
rect 19981 4536 19993 4539
rect 16209 4499 16267 4505
rect 19812 4508 19993 4536
rect 16758 4468 16764 4480
rect 15856 4440 16764 4468
rect 16758 4428 16764 4440
rect 16816 4428 16822 4480
rect 19812 4477 19840 4508
rect 19981 4505 19993 4508
rect 20027 4536 20039 4539
rect 20070 4536 20076 4548
rect 20027 4508 20076 4536
rect 20027 4505 20039 4508
rect 19981 4499 20039 4505
rect 20070 4496 20076 4508
rect 20128 4496 20134 4548
rect 20197 4539 20255 4545
rect 20197 4505 20209 4539
rect 20243 4536 20255 4539
rect 20530 4536 20536 4548
rect 20243 4508 20536 4536
rect 20243 4505 20255 4508
rect 20197 4499 20255 4505
rect 20530 4496 20536 4508
rect 20588 4496 20594 4548
rect 22796 4508 23244 4536
rect 22744 4490 22796 4496
rect 19797 4471 19855 4477
rect 19797 4437 19809 4471
rect 19843 4437 19855 4471
rect 23216 4468 23244 4508
rect 23290 4496 23296 4548
rect 23348 4496 23354 4548
rect 23477 4539 23535 4545
rect 23477 4505 23489 4539
rect 23523 4536 23535 4539
rect 24486 4536 24492 4548
rect 23523 4508 24492 4536
rect 23523 4505 23535 4508
rect 23477 4499 23535 4505
rect 23492 4468 23520 4499
rect 24486 4496 24492 4508
rect 24544 4496 24550 4548
rect 23216 4440 23520 4468
rect 24596 4468 24624 4567
rect 24688 4548 24716 4578
rect 24765 4573 24777 4578
rect 24811 4573 24823 4607
rect 24765 4567 24823 4573
rect 24854 4564 24860 4616
rect 24912 4564 24918 4616
rect 25148 4613 25176 4644
rect 25332 4644 25412 4672
rect 25332 4613 25360 4644
rect 25406 4632 25412 4644
rect 25464 4632 25470 4684
rect 26605 4675 26663 4681
rect 26605 4672 26617 4675
rect 26160 4644 26617 4672
rect 25041 4607 25099 4613
rect 25041 4573 25053 4607
rect 25087 4573 25099 4607
rect 25041 4567 25099 4573
rect 25133 4607 25191 4613
rect 25133 4573 25145 4607
rect 25179 4573 25191 4607
rect 25133 4567 25191 4573
rect 25317 4607 25375 4613
rect 25317 4573 25329 4607
rect 25363 4573 25375 4607
rect 25317 4567 25375 4573
rect 24670 4496 24676 4548
rect 24728 4496 24734 4548
rect 25056 4536 25084 4567
rect 25590 4564 25596 4616
rect 25648 4564 25654 4616
rect 26160 4613 26188 4644
rect 26605 4641 26617 4644
rect 26651 4641 26663 4675
rect 26605 4635 26663 4641
rect 26970 4632 26976 4684
rect 27028 4672 27034 4684
rect 27065 4675 27123 4681
rect 27065 4672 27077 4675
rect 27028 4644 27077 4672
rect 27028 4632 27034 4644
rect 27065 4641 27077 4644
rect 27111 4672 27123 4675
rect 27111 4644 27384 4672
rect 27111 4641 27123 4644
rect 27065 4635 27123 4641
rect 26145 4607 26203 4613
rect 26145 4573 26157 4607
rect 26191 4573 26203 4607
rect 26145 4567 26203 4573
rect 24964 4508 25084 4536
rect 25501 4539 25559 4545
rect 24964 4468 24992 4508
rect 25501 4505 25513 4539
rect 25547 4536 25559 4539
rect 26160 4536 26188 4567
rect 26326 4564 26332 4616
rect 26384 4604 26390 4616
rect 27356 4613 27384 4644
rect 27982 4632 27988 4684
rect 28040 4632 28046 4684
rect 28074 4632 28080 4684
rect 28132 4672 28138 4684
rect 28629 4675 28687 4681
rect 28629 4672 28641 4675
rect 28132 4644 28641 4672
rect 28132 4632 28138 4644
rect 28629 4641 28641 4644
rect 28675 4641 28687 4675
rect 28629 4635 28687 4641
rect 29270 4632 29276 4684
rect 29328 4632 29334 4684
rect 26697 4607 26755 4613
rect 26697 4604 26709 4607
rect 26384 4576 26709 4604
rect 26384 4564 26390 4576
rect 26697 4573 26709 4576
rect 26743 4573 26755 4607
rect 26697 4567 26755 4573
rect 27341 4607 27399 4613
rect 27341 4573 27353 4607
rect 27387 4604 27399 4607
rect 27893 4607 27951 4613
rect 27893 4604 27905 4607
rect 27387 4576 27905 4604
rect 27387 4573 27399 4576
rect 27341 4567 27399 4573
rect 27893 4573 27905 4576
rect 27939 4573 27951 4607
rect 29288 4604 29316 4632
rect 29549 4607 29607 4613
rect 29549 4604 29561 4607
rect 29288 4576 29561 4604
rect 27893 4567 27951 4573
rect 29549 4573 29561 4576
rect 29595 4573 29607 4607
rect 29549 4567 29607 4573
rect 29638 4564 29644 4616
rect 29696 4604 29702 4616
rect 30101 4607 30159 4613
rect 30101 4604 30113 4607
rect 29696 4576 30113 4604
rect 29696 4564 29702 4576
rect 30101 4573 30113 4576
rect 30147 4573 30159 4607
rect 30101 4567 30159 4573
rect 25547 4508 26188 4536
rect 26237 4539 26295 4545
rect 25547 4505 25559 4508
rect 25501 4499 25559 4505
rect 26237 4505 26249 4539
rect 26283 4536 26295 4539
rect 27157 4539 27215 4545
rect 27157 4536 27169 4539
rect 26283 4508 27169 4536
rect 26283 4505 26295 4508
rect 26237 4499 26295 4505
rect 27157 4505 27169 4508
rect 27203 4505 27215 4539
rect 30116 4536 30144 4567
rect 30282 4564 30288 4616
rect 30340 4564 30346 4616
rect 31754 4536 31760 4548
rect 30116 4508 31760 4536
rect 27157 4499 27215 4505
rect 31754 4496 31760 4508
rect 31812 4496 31818 4548
rect 24596 4440 24992 4468
rect 26421 4471 26479 4477
rect 19797 4431 19855 4437
rect 26421 4437 26433 4471
rect 26467 4468 26479 4471
rect 27706 4468 27712 4480
rect 26467 4440 27712 4468
rect 26467 4437 26479 4440
rect 26421 4431 26479 4437
rect 27706 4428 27712 4440
rect 27764 4468 27770 4480
rect 31938 4468 31944 4480
rect 27764 4440 31944 4468
rect 27764 4428 27770 4440
rect 31938 4428 31944 4440
rect 31996 4428 32002 4480
rect 1104 4378 38272 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38272 4378
rect 1104 4304 38272 4326
rect 9122 4264 9128 4276
rect 8312 4236 9128 4264
rect 8312 4205 8340 4236
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 9769 4267 9827 4273
rect 9769 4264 9781 4267
rect 9732 4236 9781 4264
rect 9732 4224 9738 4236
rect 9769 4233 9781 4236
rect 9815 4233 9827 4267
rect 9769 4227 9827 4233
rect 14458 4224 14464 4276
rect 14516 4264 14522 4276
rect 14553 4267 14611 4273
rect 14553 4264 14565 4267
rect 14516 4236 14565 4264
rect 14516 4224 14522 4236
rect 14553 4233 14565 4236
rect 14599 4233 14611 4267
rect 14553 4227 14611 4233
rect 25498 4224 25504 4276
rect 25556 4224 25562 4276
rect 27893 4267 27951 4273
rect 27893 4233 27905 4267
rect 27939 4264 27951 4267
rect 27982 4264 27988 4276
rect 27939 4236 27988 4264
rect 27939 4233 27951 4236
rect 27893 4227 27951 4233
rect 27982 4224 27988 4236
rect 28040 4224 28046 4276
rect 8297 4199 8355 4205
rect 8297 4165 8309 4199
rect 8343 4165 8355 4199
rect 8297 4159 8355 4165
rect 8570 4156 8576 4208
rect 8628 4196 8634 4208
rect 25516 4196 25544 4224
rect 8628 4168 8786 4196
rect 24964 4168 25544 4196
rect 8628 4156 8634 4168
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 8021 4131 8079 4137
rect 8021 4128 8033 4131
rect 6972 4100 8033 4128
rect 6972 4088 6978 4100
rect 8021 4097 8033 4100
rect 8067 4097 8079 4131
rect 8021 4091 8079 4097
rect 14366 4088 14372 4140
rect 14424 4088 14430 4140
rect 24964 4137 24992 4168
rect 24949 4131 25007 4137
rect 24949 4097 24961 4131
rect 24995 4097 25007 4131
rect 24949 4091 25007 4097
rect 25130 4088 25136 4140
rect 25188 4088 25194 4140
rect 25222 4088 25228 4140
rect 25280 4088 25286 4140
rect 25409 4131 25467 4137
rect 25409 4097 25421 4131
rect 25455 4128 25467 4131
rect 25516 4128 25544 4168
rect 25455 4100 25544 4128
rect 27801 4131 27859 4137
rect 25455 4097 25467 4100
rect 25409 4091 25467 4097
rect 27801 4097 27813 4131
rect 27847 4097 27859 4131
rect 27801 4091 27859 4097
rect 25317 4063 25375 4069
rect 25317 4029 25329 4063
rect 25363 4060 25375 4063
rect 26326 4060 26332 4072
rect 25363 4032 26332 4060
rect 25363 4029 25375 4032
rect 25317 4023 25375 4029
rect 26326 4020 26332 4032
rect 26384 4020 26390 4072
rect 27816 4060 27844 4091
rect 27890 4088 27896 4140
rect 27948 4128 27954 4140
rect 27985 4131 28043 4137
rect 27985 4128 27997 4131
rect 27948 4100 27997 4128
rect 27948 4088 27954 4100
rect 27985 4097 27997 4100
rect 28031 4097 28043 4131
rect 27985 4091 28043 4097
rect 30098 4088 30104 4140
rect 30156 4088 30162 4140
rect 30116 4060 30144 4088
rect 27816 4032 30144 4060
rect 25133 3995 25191 4001
rect 25133 3961 25145 3995
rect 25179 3992 25191 3995
rect 25406 3992 25412 4004
rect 25179 3964 25412 3992
rect 25179 3961 25191 3964
rect 25133 3955 25191 3961
rect 25406 3952 25412 3964
rect 25464 3992 25470 4004
rect 27816 3992 27844 4032
rect 25464 3964 27844 3992
rect 25464 3952 25470 3964
rect 1104 3834 38272 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38272 3834
rect 1104 3760 38272 3782
rect 1104 3290 38272 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38272 3290
rect 1104 3216 38272 3238
rect 17218 3136 17224 3188
rect 17276 3136 17282 3188
rect 1946 3000 1952 3052
rect 2004 3000 2010 3052
rect 2406 3000 2412 3052
rect 2464 3000 2470 3052
rect 12526 3000 12532 3052
rect 12584 3000 12590 3052
rect 13170 3000 13176 3052
rect 13228 3000 13234 3052
rect 15102 3000 15108 3052
rect 15160 3000 15166 3052
rect 17236 3049 17264 3136
rect 37550 3068 37556 3120
rect 37608 3068 37614 3120
rect 17221 3043 17279 3049
rect 17221 3009 17233 3043
rect 17267 3009 17279 3043
rect 17221 3003 17279 3009
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3040 20039 3043
rect 25958 3040 25964 3052
rect 20027 3012 25964 3040
rect 20027 3009 20039 3012
rect 19981 3003 20039 3009
rect 25958 3000 25964 3012
rect 26016 3000 26022 3052
rect 1762 2796 1768 2848
rect 1820 2796 1826 2848
rect 2222 2796 2228 2848
rect 2280 2796 2286 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 12345 2839 12403 2845
rect 12345 2836 12357 2839
rect 8444 2808 12357 2836
rect 8444 2796 8450 2808
rect 12345 2805 12357 2808
rect 12391 2805 12403 2839
rect 12345 2799 12403 2805
rect 12986 2796 12992 2848
rect 13044 2796 13050 2848
rect 14918 2796 14924 2848
rect 14976 2796 14982 2848
rect 17402 2796 17408 2848
rect 17460 2796 17466 2848
rect 19794 2796 19800 2848
rect 19852 2796 19858 2848
rect 37182 2796 37188 2848
rect 37240 2836 37246 2848
rect 37645 2839 37703 2845
rect 37645 2836 37657 2839
rect 37240 2808 37657 2836
rect 37240 2796 37246 2808
rect 37645 2805 37657 2808
rect 37691 2805 37703 2839
rect 37645 2799 37703 2805
rect 1104 2746 38272 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38272 2746
rect 1104 2672 38272 2694
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 8754 2632 8760 2644
rect 8711 2604 8760 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 10192 2604 11161 2632
rect 10192 2592 10198 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 11149 2595 11207 2601
rect 37645 2567 37703 2573
rect 37645 2564 37657 2567
rect 26206 2536 37657 2564
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 26206 2496 26234 2536
rect 37645 2533 37657 2536
rect 37691 2533 37703 2567
rect 37645 2527 37703 2533
rect 8996 2468 26234 2496
rect 8996 2456 9002 2468
rect 1762 2388 1768 2440
rect 1820 2388 1826 2440
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 2280 2400 2421 2428
rect 2280 2388 2286 2400
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4798 2428 4804 2440
rect 4387 2400 4804 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 8386 2428 8392 2440
rect 6963 2400 8392 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 12986 2388 12992 2440
rect 13044 2428 13050 2440
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 13044 2400 13093 2428
rect 13044 2388 13050 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 15013 2431 15071 2437
rect 15013 2428 15025 2431
rect 14976 2400 15025 2428
rect 14976 2388 14982 2400
rect 15013 2397 15025 2400
rect 15059 2397 15071 2431
rect 15013 2391 15071 2397
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 17460 2400 17601 2428
rect 17460 2388 17466 2400
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 19794 2388 19800 2440
rect 19852 2388 19858 2440
rect 37458 2388 37464 2440
rect 37516 2388 37522 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 72 2332 1409 2360
rect 72 2320 78 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 2038 2320 2044 2372
rect 2096 2320 2102 2372
rect 3970 2320 3976 2372
rect 4028 2320 4034 2372
rect 6546 2320 6552 2372
rect 6604 2320 6610 2372
rect 10962 2320 10968 2372
rect 11020 2360 11026 2372
rect 11241 2363 11299 2369
rect 11241 2360 11253 2363
rect 11020 2332 11253 2360
rect 11020 2320 11026 2332
rect 11241 2329 11253 2332
rect 11287 2329 11299 2363
rect 11241 2323 11299 2329
rect 14642 2320 14648 2372
rect 14700 2360 14706 2372
rect 14700 2332 19380 2360
rect 14700 2320 14706 2332
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 15010 2252 15016 2304
rect 15068 2292 15074 2304
rect 15289 2295 15347 2301
rect 15289 2292 15301 2295
rect 15068 2264 15301 2292
rect 15068 2252 15074 2264
rect 15289 2261 15301 2264
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 19352 2292 19380 2332
rect 19426 2320 19432 2372
rect 19484 2320 19490 2372
rect 27065 2363 27123 2369
rect 27065 2360 27077 2363
rect 26206 2332 27077 2360
rect 26206 2292 26234 2332
rect 27065 2329 27077 2332
rect 27111 2329 27123 2363
rect 27065 2323 27123 2329
rect 19352 2264 26234 2292
rect 17681 2255 17739 2261
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26476 2264 27169 2292
rect 26476 2252 26482 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 1104 2202 38272 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38272 2202
rect 1104 2128 38272 2150
<< via1 >>
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 20 39040 72 39092
rect 4896 39083 4948 39092
rect 4896 39049 4905 39083
rect 4905 39049 4939 39083
rect 4939 39049 4948 39083
rect 4896 39040 4948 39049
rect 9036 39040 9088 39092
rect 11060 39040 11112 39092
rect 13176 39083 13228 39092
rect 13176 39049 13185 39083
rect 13185 39049 13219 39083
rect 13219 39049 13228 39083
rect 13176 39040 13228 39049
rect 17408 39040 17460 39092
rect 21916 39040 21968 39092
rect 26424 39040 26476 39092
rect 33140 39083 33192 39092
rect 33140 39049 33149 39083
rect 33149 39049 33183 39083
rect 33183 39049 33192 39083
rect 33140 39040 33192 39049
rect 35440 39040 35492 39092
rect 12348 38972 12400 39024
rect 15476 38972 15528 39024
rect 30932 38972 30984 39024
rect 1768 38947 1820 38956
rect 1768 38913 1777 38947
rect 1777 38913 1811 38947
rect 1811 38913 1820 38947
rect 1768 38904 1820 38913
rect 5080 38947 5132 38956
rect 5080 38913 5089 38947
rect 5089 38913 5123 38947
rect 5123 38913 5132 38947
rect 5080 38904 5132 38913
rect 9220 38947 9272 38956
rect 9220 38913 9229 38947
rect 9229 38913 9263 38947
rect 9263 38913 9272 38947
rect 9220 38904 9272 38913
rect 12072 38947 12124 38956
rect 12072 38913 12081 38947
rect 12081 38913 12115 38947
rect 12115 38913 12124 38947
rect 12072 38904 12124 38913
rect 12440 38904 12492 38956
rect 17960 38947 18012 38956
rect 17960 38913 17969 38947
rect 17969 38913 18003 38947
rect 18003 38913 18012 38947
rect 17960 38904 18012 38913
rect 19432 38947 19484 38956
rect 19432 38913 19441 38947
rect 19441 38913 19475 38947
rect 19475 38913 19484 38947
rect 19432 38904 19484 38913
rect 20076 38947 20128 38956
rect 20076 38913 20085 38947
rect 20085 38913 20119 38947
rect 20119 38913 20128 38947
rect 20076 38904 20128 38913
rect 22376 38947 22428 38956
rect 22376 38913 22385 38947
rect 22385 38913 22419 38947
rect 22419 38913 22428 38947
rect 22376 38904 22428 38913
rect 27068 38947 27120 38956
rect 27068 38913 27077 38947
rect 27077 38913 27111 38947
rect 27111 38913 27120 38947
rect 27068 38904 27120 38913
rect 27712 38947 27764 38956
rect 27712 38913 27721 38947
rect 27721 38913 27755 38947
rect 27755 38913 27764 38947
rect 27712 38904 27764 38913
rect 33048 38947 33100 38956
rect 33048 38913 33057 38947
rect 33057 38913 33091 38947
rect 33091 38913 33100 38947
rect 33048 38904 33100 38913
rect 35624 38947 35676 38956
rect 35624 38913 35633 38947
rect 35633 38913 35667 38947
rect 35667 38913 35676 38947
rect 35624 38904 35676 38913
rect 37372 38904 37424 38956
rect 20352 38879 20404 38888
rect 20352 38845 20361 38879
rect 20361 38845 20395 38879
rect 20395 38845 20404 38879
rect 20352 38836 20404 38845
rect 15568 38811 15620 38820
rect 15568 38777 15577 38811
rect 15577 38777 15611 38811
rect 15611 38777 15620 38811
rect 15568 38768 15620 38777
rect 29736 38768 29788 38820
rect 37648 38811 37700 38820
rect 37648 38777 37657 38811
rect 37657 38777 37691 38811
rect 37691 38777 37700 38811
rect 37648 38768 37700 38777
rect 12808 38700 12860 38752
rect 19616 38743 19668 38752
rect 19616 38709 19625 38743
rect 19625 38709 19659 38743
rect 19659 38709 19668 38743
rect 19616 38700 19668 38709
rect 27620 38743 27672 38752
rect 27620 38709 27629 38743
rect 27629 38709 27663 38743
rect 27663 38709 27672 38743
rect 27620 38700 27672 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 5080 38496 5132 38548
rect 9220 38496 9272 38548
rect 17960 38496 18012 38548
rect 5172 38335 5224 38344
rect 5172 38301 5181 38335
rect 5181 38301 5215 38335
rect 5215 38301 5224 38335
rect 5172 38292 5224 38301
rect 8576 38335 8628 38344
rect 8576 38301 8585 38335
rect 8585 38301 8619 38335
rect 8619 38301 8628 38335
rect 8576 38292 8628 38301
rect 9036 38335 9088 38344
rect 9036 38301 9045 38335
rect 9045 38301 9079 38335
rect 9079 38301 9088 38335
rect 9036 38292 9088 38301
rect 11336 38292 11388 38344
rect 13728 38292 13780 38344
rect 19616 38360 19668 38412
rect 24860 38360 24912 38412
rect 9588 38267 9640 38276
rect 9588 38233 9597 38267
rect 9597 38233 9631 38267
rect 9631 38233 9640 38267
rect 9588 38224 9640 38233
rect 10232 38224 10284 38276
rect 11060 38224 11112 38276
rect 12808 38267 12860 38276
rect 12808 38233 12817 38267
rect 12817 38233 12851 38267
rect 12851 38233 12860 38267
rect 12808 38224 12860 38233
rect 12900 38224 12952 38276
rect 20812 38292 20864 38344
rect 21272 38335 21324 38344
rect 21272 38301 21281 38335
rect 21281 38301 21315 38335
rect 21315 38301 21324 38335
rect 21272 38292 21324 38301
rect 27712 38496 27764 38548
rect 26056 38360 26108 38412
rect 11888 38156 11940 38208
rect 13728 38156 13780 38208
rect 20996 38199 21048 38208
rect 20996 38165 21005 38199
rect 21005 38165 21039 38199
rect 21039 38165 21048 38199
rect 20996 38156 21048 38165
rect 22008 38156 22060 38208
rect 24032 38156 24084 38208
rect 25596 38267 25648 38276
rect 25596 38233 25605 38267
rect 25605 38233 25639 38267
rect 25639 38233 25648 38267
rect 25596 38224 25648 38233
rect 26056 38224 26108 38276
rect 26976 38156 27028 38208
rect 27620 38360 27672 38412
rect 33048 38496 33100 38548
rect 35624 38496 35676 38548
rect 37924 38496 37976 38548
rect 32680 38360 32732 38412
rect 29552 38335 29604 38344
rect 29552 38301 29561 38335
rect 29561 38301 29595 38335
rect 29595 38301 29604 38335
rect 29552 38292 29604 38301
rect 29644 38335 29696 38344
rect 29644 38301 29653 38335
rect 29653 38301 29687 38335
rect 29687 38301 29696 38335
rect 29644 38292 29696 38301
rect 31668 38292 31720 38344
rect 27528 38267 27580 38276
rect 27528 38233 27537 38267
rect 27537 38233 27571 38267
rect 27571 38233 27580 38267
rect 27528 38224 27580 38233
rect 29276 38267 29328 38276
rect 29276 38233 29285 38267
rect 29285 38233 29319 38267
rect 29319 38233 29328 38267
rect 29276 38224 29328 38233
rect 29460 38224 29512 38276
rect 28540 38156 28592 38208
rect 30380 38156 30432 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 9588 37952 9640 38004
rect 12072 37952 12124 38004
rect 12348 37995 12400 38004
rect 12348 37961 12357 37995
rect 12357 37961 12391 37995
rect 12391 37961 12400 37995
rect 12348 37952 12400 37961
rect 10692 37927 10744 37936
rect 10692 37893 10701 37927
rect 10701 37893 10735 37927
rect 10735 37893 10744 37927
rect 10692 37884 10744 37893
rect 11888 37927 11940 37936
rect 11888 37893 11897 37927
rect 11897 37893 11931 37927
rect 11931 37893 11940 37927
rect 11888 37884 11940 37893
rect 11336 37816 11388 37868
rect 12532 37859 12584 37868
rect 12532 37825 12541 37859
rect 12541 37825 12575 37859
rect 12575 37825 12584 37859
rect 12532 37816 12584 37825
rect 10784 37791 10836 37800
rect 10784 37757 10793 37791
rect 10793 37757 10827 37791
rect 10827 37757 10836 37791
rect 10784 37748 10836 37757
rect 11704 37791 11756 37800
rect 11704 37757 11713 37791
rect 11713 37757 11747 37791
rect 11747 37757 11756 37791
rect 11704 37748 11756 37757
rect 13268 37859 13320 37868
rect 13268 37825 13277 37859
rect 13277 37825 13311 37859
rect 13311 37825 13320 37859
rect 13268 37816 13320 37825
rect 15292 37952 15344 38004
rect 16304 37952 16356 38004
rect 14280 37884 14332 37936
rect 13820 37859 13872 37868
rect 13820 37825 13829 37859
rect 13829 37825 13863 37859
rect 13863 37825 13872 37859
rect 13820 37816 13872 37825
rect 14372 37859 14424 37868
rect 14372 37825 14376 37859
rect 14376 37825 14410 37859
rect 14410 37825 14424 37859
rect 14372 37816 14424 37825
rect 14556 37859 14608 37868
rect 14556 37825 14565 37859
rect 14565 37825 14599 37859
rect 14599 37825 14608 37859
rect 14556 37816 14608 37825
rect 14096 37680 14148 37732
rect 16028 37816 16080 37868
rect 16120 37859 16172 37868
rect 16120 37825 16129 37859
rect 16129 37825 16163 37859
rect 16163 37825 16172 37859
rect 16120 37816 16172 37825
rect 16212 37859 16264 37868
rect 16212 37825 16221 37859
rect 16221 37825 16255 37859
rect 16255 37825 16264 37859
rect 16212 37816 16264 37825
rect 16488 37816 16540 37868
rect 19432 37995 19484 38004
rect 19432 37961 19441 37995
rect 19441 37961 19475 37995
rect 19475 37961 19484 37995
rect 19432 37952 19484 37961
rect 20996 37952 21048 38004
rect 21272 37952 21324 38004
rect 22468 37995 22520 38004
rect 22468 37961 22477 37995
rect 22477 37961 22511 37995
rect 22511 37961 22520 37995
rect 22468 37952 22520 37961
rect 22744 37952 22796 38004
rect 24860 37995 24912 38004
rect 24860 37961 24869 37995
rect 24869 37961 24903 37995
rect 24903 37961 24912 37995
rect 24860 37952 24912 37961
rect 25596 37952 25648 38004
rect 27528 37952 27580 38004
rect 29460 37952 29512 38004
rect 29644 37952 29696 38004
rect 16856 37859 16908 37868
rect 16856 37825 16865 37859
rect 16865 37825 16899 37859
rect 16899 37825 16908 37859
rect 16856 37816 16908 37825
rect 17224 37859 17276 37868
rect 17224 37825 17233 37859
rect 17233 37825 17267 37859
rect 17267 37825 17276 37859
rect 17224 37816 17276 37825
rect 17684 37816 17736 37868
rect 17868 37816 17920 37868
rect 20812 37816 20864 37868
rect 22008 37816 22060 37868
rect 12808 37612 12860 37664
rect 16488 37655 16540 37664
rect 16488 37621 16497 37655
rect 16497 37621 16531 37655
rect 16531 37621 16540 37655
rect 16488 37612 16540 37621
rect 17960 37612 18012 37664
rect 19984 37748 20036 37800
rect 20444 37748 20496 37800
rect 22652 37791 22704 37800
rect 19294 37680 19346 37732
rect 22652 37757 22661 37791
rect 22661 37757 22695 37791
rect 22695 37757 22704 37791
rect 22652 37748 22704 37757
rect 20720 37680 20772 37732
rect 22468 37680 22520 37732
rect 25780 37927 25832 37936
rect 25780 37893 25789 37927
rect 25789 37893 25823 37927
rect 25823 37893 25832 37927
rect 25780 37884 25832 37893
rect 23112 37816 23164 37868
rect 23664 37859 23716 37868
rect 23664 37825 23673 37859
rect 23673 37825 23707 37859
rect 23707 37825 23716 37859
rect 23664 37816 23716 37825
rect 23756 37859 23808 37868
rect 23756 37825 23765 37859
rect 23765 37825 23799 37859
rect 23799 37825 23808 37859
rect 23756 37816 23808 37825
rect 25320 37859 25372 37868
rect 25320 37825 25329 37859
rect 25329 37825 25363 37859
rect 25363 37825 25372 37859
rect 25320 37816 25372 37825
rect 25228 37791 25280 37800
rect 25228 37757 25237 37791
rect 25237 37757 25271 37791
rect 25271 37757 25280 37791
rect 25228 37748 25280 37757
rect 26424 37859 26476 37868
rect 26424 37825 26433 37859
rect 26433 37825 26467 37859
rect 26467 37825 26476 37859
rect 26424 37816 26476 37825
rect 26608 37859 26660 37868
rect 26608 37825 26617 37859
rect 26617 37825 26651 37859
rect 26651 37825 26660 37859
rect 26608 37816 26660 37825
rect 29000 37816 29052 37868
rect 30380 37884 30432 37936
rect 31208 37859 31260 37868
rect 31208 37825 31217 37859
rect 31217 37825 31251 37859
rect 31251 37825 31260 37859
rect 31208 37816 31260 37825
rect 25596 37748 25648 37800
rect 26148 37791 26200 37800
rect 26148 37757 26157 37791
rect 26157 37757 26191 37791
rect 26191 37757 26200 37791
rect 26148 37748 26200 37757
rect 27068 37748 27120 37800
rect 27988 37791 28040 37800
rect 27988 37757 27997 37791
rect 27997 37757 28031 37791
rect 28031 37757 28040 37791
rect 27988 37748 28040 37757
rect 29460 37748 29512 37800
rect 31668 37748 31720 37800
rect 22376 37612 22428 37664
rect 23940 37655 23992 37664
rect 23940 37621 23949 37655
rect 23949 37621 23983 37655
rect 23983 37621 23992 37655
rect 23940 37612 23992 37621
rect 24032 37612 24084 37664
rect 25688 37612 25740 37664
rect 30932 37612 30984 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 9588 37408 9640 37460
rect 11060 37408 11112 37460
rect 16488 37408 16540 37460
rect 17868 37408 17920 37460
rect 22376 37408 22428 37460
rect 9588 37272 9640 37324
rect 15844 37272 15896 37324
rect 16028 37272 16080 37324
rect 8300 37247 8352 37256
rect 8300 37213 8309 37247
rect 8309 37213 8343 37247
rect 8343 37213 8352 37247
rect 8300 37204 8352 37213
rect 940 37136 992 37188
rect 7196 37136 7248 37188
rect 10232 37204 10284 37256
rect 17868 37315 17920 37324
rect 17868 37281 17877 37315
rect 17877 37281 17911 37315
rect 17911 37281 17920 37315
rect 17868 37272 17920 37281
rect 24860 37340 24912 37392
rect 26424 37408 26476 37460
rect 26608 37408 26660 37460
rect 22928 37315 22980 37324
rect 22928 37281 22937 37315
rect 22937 37281 22971 37315
rect 22971 37281 22980 37315
rect 22928 37272 22980 37281
rect 23480 37272 23532 37324
rect 18420 37204 18472 37256
rect 17776 37179 17828 37188
rect 17776 37145 17785 37179
rect 17785 37145 17819 37179
rect 17819 37145 17828 37179
rect 17776 37136 17828 37145
rect 20168 37247 20220 37256
rect 20168 37213 20177 37247
rect 20177 37213 20211 37247
rect 20211 37213 20220 37247
rect 20168 37204 20220 37213
rect 22744 37247 22796 37256
rect 22744 37213 22753 37247
rect 22753 37213 22787 37247
rect 22787 37213 22796 37247
rect 22744 37204 22796 37213
rect 23296 37247 23348 37256
rect 23296 37213 23305 37247
rect 23305 37213 23339 37247
rect 23339 37213 23348 37247
rect 23296 37204 23348 37213
rect 24400 37204 24452 37256
rect 27896 37272 27948 37324
rect 28632 37272 28684 37324
rect 29552 37272 29604 37324
rect 10600 37068 10652 37120
rect 17132 37068 17184 37120
rect 20720 37179 20772 37188
rect 20720 37145 20729 37179
rect 20729 37145 20763 37179
rect 20763 37145 20772 37179
rect 20720 37136 20772 37145
rect 22008 37136 22060 37188
rect 22836 37179 22888 37188
rect 18512 37068 18564 37120
rect 22836 37145 22845 37179
rect 22845 37145 22879 37179
rect 22879 37145 22888 37179
rect 22836 37136 22888 37145
rect 22376 37111 22428 37120
rect 22376 37077 22385 37111
rect 22385 37077 22419 37111
rect 22419 37077 22428 37111
rect 22376 37068 22428 37077
rect 23572 37179 23624 37188
rect 23572 37145 23581 37179
rect 23581 37145 23615 37179
rect 23615 37145 23624 37179
rect 23572 37136 23624 37145
rect 24676 37136 24728 37188
rect 27344 37204 27396 37256
rect 29276 37204 29328 37256
rect 30932 37272 30984 37324
rect 32588 37247 32640 37256
rect 32588 37213 32597 37247
rect 32597 37213 32631 37247
rect 32631 37213 32640 37247
rect 32588 37204 32640 37213
rect 26976 37136 27028 37188
rect 27988 37136 28040 37188
rect 30472 37136 30524 37188
rect 31484 37136 31536 37188
rect 24584 37068 24636 37120
rect 27620 37068 27672 37120
rect 30012 37068 30064 37120
rect 32496 37111 32548 37120
rect 32496 37077 32505 37111
rect 32505 37077 32539 37111
rect 32539 37077 32548 37111
rect 32496 37068 32548 37077
rect 37832 37111 37884 37120
rect 37832 37077 37841 37111
rect 37841 37077 37875 37111
rect 37875 37077 37884 37111
rect 37832 37068 37884 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 8300 36864 8352 36916
rect 10692 36864 10744 36916
rect 20720 36864 20772 36916
rect 9588 36796 9640 36848
rect 10600 36796 10652 36848
rect 14280 36728 14332 36780
rect 14832 36728 14884 36780
rect 17500 36728 17552 36780
rect 18420 36728 18472 36780
rect 19984 36728 20036 36780
rect 22376 36864 22428 36916
rect 22468 36728 22520 36780
rect 23480 36728 23532 36780
rect 9496 36660 9548 36712
rect 9864 36703 9916 36712
rect 9864 36669 9873 36703
rect 9873 36669 9907 36703
rect 9907 36669 9916 36703
rect 9864 36660 9916 36669
rect 17040 36660 17092 36712
rect 19156 36660 19208 36712
rect 20720 36660 20772 36712
rect 25136 36864 25188 36916
rect 27804 36864 27856 36916
rect 29000 36864 29052 36916
rect 30012 36864 30064 36916
rect 31208 36864 31260 36916
rect 31484 36864 31536 36916
rect 32496 36864 32548 36916
rect 23940 36728 23992 36780
rect 24492 36771 24544 36780
rect 24492 36737 24501 36771
rect 24501 36737 24535 36771
rect 24535 36737 24544 36771
rect 24492 36728 24544 36737
rect 27712 36771 27764 36780
rect 27712 36737 27721 36771
rect 27721 36737 27755 36771
rect 27755 36737 27764 36771
rect 27712 36728 27764 36737
rect 22560 36592 22612 36644
rect 23480 36592 23532 36644
rect 27896 36660 27948 36712
rect 28264 36771 28316 36780
rect 28264 36737 28273 36771
rect 28273 36737 28307 36771
rect 28307 36737 28316 36771
rect 28264 36728 28316 36737
rect 29368 36728 29420 36780
rect 28172 36660 28224 36712
rect 29460 36660 29512 36712
rect 29644 36703 29696 36712
rect 29644 36669 29653 36703
rect 29653 36669 29687 36703
rect 29687 36669 29696 36703
rect 29644 36660 29696 36669
rect 23940 36592 23992 36644
rect 24124 36592 24176 36644
rect 7472 36524 7524 36576
rect 11520 36524 11572 36576
rect 15660 36524 15712 36576
rect 15752 36524 15804 36576
rect 17960 36524 18012 36576
rect 25136 36592 25188 36644
rect 29276 36592 29328 36644
rect 24584 36567 24636 36576
rect 24584 36533 24593 36567
rect 24593 36533 24627 36567
rect 24627 36533 24636 36567
rect 24584 36524 24636 36533
rect 26240 36524 26292 36576
rect 27436 36524 27488 36576
rect 28448 36567 28500 36576
rect 28448 36533 28457 36567
rect 28457 36533 28491 36567
rect 28491 36533 28500 36567
rect 28448 36524 28500 36533
rect 28632 36524 28684 36576
rect 30656 36703 30708 36712
rect 30656 36669 30665 36703
rect 30665 36669 30699 36703
rect 30699 36669 30708 36703
rect 30656 36660 30708 36669
rect 33692 36728 33744 36780
rect 32220 36660 32272 36712
rect 33140 36524 33192 36576
rect 34060 36567 34112 36576
rect 34060 36533 34069 36567
rect 34069 36533 34103 36567
rect 34103 36533 34112 36567
rect 34060 36524 34112 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 13176 36320 13228 36372
rect 13636 36320 13688 36372
rect 13820 36320 13872 36372
rect 14556 36320 14608 36372
rect 15200 36320 15252 36372
rect 15292 36363 15344 36372
rect 15292 36329 15301 36363
rect 15301 36329 15335 36363
rect 15335 36329 15344 36363
rect 15292 36320 15344 36329
rect 16764 36320 16816 36372
rect 17776 36320 17828 36372
rect 11704 36252 11756 36304
rect 6828 36184 6880 36236
rect 7472 36184 7524 36236
rect 5724 36159 5776 36168
rect 5724 36125 5733 36159
rect 5733 36125 5767 36159
rect 5767 36125 5776 36159
rect 5724 36116 5776 36125
rect 6276 36091 6328 36100
rect 6276 36057 6285 36091
rect 6285 36057 6319 36091
rect 6319 36057 6328 36091
rect 6276 36048 6328 36057
rect 9036 36116 9088 36168
rect 9772 36159 9824 36168
rect 9772 36125 9781 36159
rect 9781 36125 9815 36159
rect 9815 36125 9824 36159
rect 9772 36116 9824 36125
rect 10232 36116 10284 36168
rect 10600 36116 10652 36168
rect 11336 36116 11388 36168
rect 11520 36159 11572 36168
rect 11520 36125 11529 36159
rect 11529 36125 11563 36159
rect 11563 36125 11572 36159
rect 11520 36116 11572 36125
rect 11888 36116 11940 36168
rect 7748 36023 7800 36032
rect 7748 35989 7757 36023
rect 7757 35989 7791 36023
rect 7791 35989 7800 36023
rect 7748 35980 7800 35989
rect 9404 36023 9456 36032
rect 9404 35989 9413 36023
rect 9413 35989 9447 36023
rect 9447 35989 9456 36023
rect 9404 35980 9456 35989
rect 9588 36023 9640 36032
rect 9588 35989 9597 36023
rect 9597 35989 9631 36023
rect 9631 35989 9640 36023
rect 9588 35980 9640 35989
rect 11796 36048 11848 36100
rect 12256 36116 12308 36168
rect 11980 35980 12032 36032
rect 12808 35980 12860 36032
rect 12992 36091 13044 36100
rect 12992 36057 13001 36091
rect 13001 36057 13035 36091
rect 13035 36057 13044 36091
rect 12992 36048 13044 36057
rect 13176 36116 13228 36168
rect 14096 36116 14148 36168
rect 14280 36159 14332 36168
rect 14280 36125 14289 36159
rect 14289 36125 14323 36159
rect 14323 36125 14332 36159
rect 14280 36116 14332 36125
rect 17132 36252 17184 36304
rect 14556 36091 14608 36100
rect 14556 36057 14565 36091
rect 14565 36057 14599 36091
rect 14599 36057 14608 36091
rect 14556 36048 14608 36057
rect 14832 36116 14884 36168
rect 15660 36159 15712 36168
rect 15660 36125 15669 36159
rect 15669 36125 15703 36159
rect 15703 36125 15712 36159
rect 15660 36116 15712 36125
rect 15752 36159 15804 36168
rect 15752 36125 15761 36159
rect 15761 36125 15795 36159
rect 15795 36125 15804 36159
rect 15752 36116 15804 36125
rect 15108 36048 15160 36100
rect 15568 36091 15620 36100
rect 15568 36057 15577 36091
rect 15577 36057 15611 36091
rect 15611 36057 15620 36091
rect 15568 36048 15620 36057
rect 16212 36159 16264 36168
rect 16212 36125 16221 36159
rect 16221 36125 16255 36159
rect 16255 36125 16264 36159
rect 16212 36116 16264 36125
rect 16672 36116 16724 36168
rect 16764 36159 16816 36168
rect 16764 36125 16773 36159
rect 16773 36125 16807 36159
rect 16807 36125 16816 36159
rect 16764 36116 16816 36125
rect 16856 36159 16908 36168
rect 16856 36125 16866 36159
rect 16866 36125 16900 36159
rect 16900 36125 16908 36159
rect 16856 36116 16908 36125
rect 17224 36159 17276 36168
rect 17960 36184 18012 36236
rect 17224 36125 17238 36159
rect 17238 36125 17272 36159
rect 17272 36125 17276 36159
rect 17224 36116 17276 36125
rect 15844 35980 15896 36032
rect 16120 36091 16172 36100
rect 16120 36057 16129 36091
rect 16129 36057 16163 36091
rect 16163 36057 16172 36091
rect 16120 36048 16172 36057
rect 17040 36091 17092 36100
rect 17040 36057 17049 36091
rect 17049 36057 17083 36091
rect 17083 36057 17092 36091
rect 17040 36048 17092 36057
rect 17132 36091 17184 36100
rect 17132 36057 17141 36091
rect 17141 36057 17175 36091
rect 17175 36057 17184 36091
rect 17132 36048 17184 36057
rect 17868 36159 17920 36168
rect 17868 36125 17877 36159
rect 17877 36125 17911 36159
rect 17911 36125 17920 36159
rect 17868 36116 17920 36125
rect 18052 36116 18104 36168
rect 22468 36320 22520 36372
rect 23020 36320 23072 36372
rect 23572 36320 23624 36372
rect 23756 36320 23808 36372
rect 24308 36320 24360 36372
rect 28264 36320 28316 36372
rect 29276 36320 29328 36372
rect 30656 36320 30708 36372
rect 32220 36363 32272 36372
rect 32220 36329 32229 36363
rect 32229 36329 32263 36363
rect 32263 36329 32272 36363
rect 32220 36320 32272 36329
rect 34060 36320 34112 36372
rect 19984 36252 20036 36304
rect 23940 36252 23992 36304
rect 24492 36252 24544 36304
rect 19340 36184 19392 36236
rect 22100 36184 22152 36236
rect 23296 36184 23348 36236
rect 30012 36252 30064 36304
rect 17592 36048 17644 36100
rect 22836 36116 22888 36168
rect 23204 36116 23256 36168
rect 24584 36116 24636 36168
rect 19064 36048 19116 36100
rect 19984 36091 20036 36100
rect 19984 36057 19993 36091
rect 19993 36057 20027 36091
rect 20027 36057 20036 36091
rect 19984 36048 20036 36057
rect 20536 36048 20588 36100
rect 21088 36048 21140 36100
rect 17408 36023 17460 36032
rect 17408 35989 17417 36023
rect 17417 35989 17451 36023
rect 17451 35989 17460 36023
rect 17408 35980 17460 35989
rect 18604 36023 18656 36032
rect 18604 35989 18613 36023
rect 18613 35989 18647 36023
rect 18647 35989 18656 36023
rect 18604 35980 18656 35989
rect 22928 35980 22980 36032
rect 24952 36048 25004 36100
rect 25964 36116 26016 36168
rect 27252 36159 27304 36168
rect 27252 36125 27261 36159
rect 27261 36125 27295 36159
rect 27295 36125 27304 36159
rect 27252 36116 27304 36125
rect 27344 36159 27396 36168
rect 27344 36125 27354 36159
rect 27354 36125 27388 36159
rect 27388 36125 27396 36159
rect 27988 36184 28040 36236
rect 28724 36227 28776 36236
rect 28724 36193 28733 36227
rect 28733 36193 28767 36227
rect 28767 36193 28776 36227
rect 28724 36184 28776 36193
rect 27344 36116 27396 36125
rect 28264 36116 28316 36168
rect 28540 36159 28592 36168
rect 28540 36125 28549 36159
rect 28549 36125 28583 36159
rect 28583 36125 28592 36159
rect 28540 36116 28592 36125
rect 26056 36023 26108 36032
rect 26056 35989 26065 36023
rect 26065 35989 26099 36023
rect 26099 35989 26108 36023
rect 26056 35980 26108 35989
rect 26424 36048 26476 36100
rect 29828 36048 29880 36100
rect 30840 36048 30892 36100
rect 30748 35980 30800 36032
rect 33140 35980 33192 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 6276 35776 6328 35828
rect 7748 35776 7800 35828
rect 8116 35776 8168 35828
rect 9128 35776 9180 35828
rect 12900 35776 12952 35828
rect 9588 35708 9640 35760
rect 10232 35708 10284 35760
rect 11152 35708 11204 35760
rect 12992 35708 13044 35760
rect 7472 35572 7524 35624
rect 8208 35572 8260 35624
rect 8300 35615 8352 35624
rect 8300 35581 8309 35615
rect 8309 35581 8343 35615
rect 8343 35581 8352 35615
rect 8300 35572 8352 35581
rect 9220 35683 9272 35692
rect 9220 35649 9229 35683
rect 9229 35649 9263 35683
rect 9263 35649 9272 35683
rect 9220 35640 9272 35649
rect 13360 35776 13412 35828
rect 14280 35776 14332 35828
rect 18604 35708 18656 35760
rect 20444 35708 20496 35760
rect 22192 35751 22244 35760
rect 22192 35717 22201 35751
rect 22201 35717 22235 35751
rect 22235 35717 22244 35751
rect 22192 35708 22244 35717
rect 13544 35683 13596 35692
rect 13544 35649 13553 35683
rect 13553 35649 13587 35683
rect 13587 35649 13596 35683
rect 13544 35640 13596 35649
rect 13728 35683 13780 35692
rect 13728 35649 13737 35683
rect 13737 35649 13771 35683
rect 13771 35649 13780 35683
rect 13728 35640 13780 35649
rect 9496 35572 9548 35624
rect 13636 35572 13688 35624
rect 18880 35683 18932 35692
rect 18880 35649 18889 35683
rect 18889 35649 18923 35683
rect 18923 35649 18932 35683
rect 18880 35640 18932 35649
rect 16212 35572 16264 35624
rect 17960 35572 18012 35624
rect 11336 35504 11388 35556
rect 19984 35640 20036 35692
rect 20076 35640 20128 35692
rect 21180 35683 21232 35692
rect 21180 35649 21189 35683
rect 21189 35649 21223 35683
rect 21223 35649 21232 35683
rect 21180 35640 21232 35649
rect 22100 35683 22152 35692
rect 22100 35649 22107 35683
rect 22107 35649 22152 35683
rect 22100 35640 22152 35649
rect 22284 35683 22336 35692
rect 22284 35649 22290 35683
rect 22290 35649 22324 35683
rect 22324 35649 22336 35683
rect 22284 35640 22336 35649
rect 22376 35683 22428 35692
rect 22376 35649 22390 35683
rect 22390 35649 22424 35683
rect 22424 35649 22428 35683
rect 22376 35640 22428 35649
rect 22560 35640 22612 35692
rect 22836 35683 22888 35692
rect 22836 35649 22845 35683
rect 22845 35649 22879 35683
rect 22879 35649 22888 35683
rect 22836 35640 22888 35649
rect 22928 35683 22980 35692
rect 22928 35649 22938 35683
rect 22938 35649 22972 35683
rect 22972 35649 22980 35683
rect 23296 35776 23348 35828
rect 23664 35776 23716 35828
rect 23204 35751 23256 35760
rect 23204 35717 23213 35751
rect 23213 35717 23247 35751
rect 23247 35717 23256 35751
rect 23204 35708 23256 35717
rect 24032 35708 24084 35760
rect 22928 35640 22980 35649
rect 21456 35572 21508 35624
rect 22744 35572 22796 35624
rect 23756 35683 23808 35692
rect 23756 35649 23765 35683
rect 23765 35649 23799 35683
rect 23799 35649 23808 35683
rect 23756 35640 23808 35649
rect 25136 35751 25188 35760
rect 25136 35717 25145 35751
rect 25145 35717 25179 35751
rect 25179 35717 25188 35751
rect 25136 35708 25188 35717
rect 23848 35572 23900 35624
rect 24860 35683 24912 35692
rect 24860 35649 24869 35683
rect 24869 35649 24903 35683
rect 24903 35649 24912 35683
rect 24860 35640 24912 35649
rect 24952 35640 25004 35692
rect 25964 35776 26016 35828
rect 26056 35776 26108 35828
rect 27804 35776 27856 35828
rect 25412 35640 25464 35692
rect 25872 35640 25924 35692
rect 28724 35708 28776 35760
rect 26056 35683 26108 35692
rect 26056 35649 26065 35683
rect 26065 35649 26099 35683
rect 26099 35649 26108 35683
rect 26056 35640 26108 35649
rect 26516 35683 26568 35692
rect 26516 35649 26525 35683
rect 26525 35649 26559 35683
rect 26559 35649 26568 35683
rect 26516 35640 26568 35649
rect 27344 35640 27396 35692
rect 30472 35708 30524 35760
rect 20996 35504 21048 35556
rect 23664 35504 23716 35556
rect 27436 35615 27488 35624
rect 27436 35581 27445 35615
rect 27445 35581 27479 35615
rect 27479 35581 27488 35615
rect 27436 35572 27488 35581
rect 28172 35572 28224 35624
rect 28264 35572 28316 35624
rect 28448 35572 28500 35624
rect 29828 35640 29880 35692
rect 30012 35683 30064 35692
rect 30012 35649 30021 35683
rect 30021 35649 30055 35683
rect 30055 35649 30064 35683
rect 30012 35640 30064 35649
rect 25872 35504 25924 35556
rect 10968 35479 11020 35488
rect 10968 35445 10977 35479
rect 10977 35445 11011 35479
rect 11011 35445 11020 35479
rect 10968 35436 11020 35445
rect 12532 35436 12584 35488
rect 18696 35479 18748 35488
rect 18696 35445 18705 35479
rect 18705 35445 18739 35479
rect 18739 35445 18748 35479
rect 18696 35436 18748 35445
rect 19340 35436 19392 35488
rect 23480 35479 23532 35488
rect 23480 35445 23489 35479
rect 23489 35445 23523 35479
rect 23523 35445 23532 35479
rect 23480 35436 23532 35445
rect 23940 35436 23992 35488
rect 25504 35479 25556 35488
rect 25504 35445 25513 35479
rect 25513 35445 25547 35479
rect 25547 35445 25556 35479
rect 25504 35436 25556 35445
rect 26608 35436 26660 35488
rect 30748 35819 30800 35828
rect 30748 35785 30757 35819
rect 30757 35785 30791 35819
rect 30791 35785 30800 35819
rect 30748 35776 30800 35785
rect 32588 35708 32640 35760
rect 31392 35683 31444 35692
rect 31392 35649 31401 35683
rect 31401 35649 31435 35683
rect 31435 35649 31444 35683
rect 31392 35640 31444 35649
rect 33508 35683 33560 35692
rect 33508 35649 33517 35683
rect 33517 35649 33551 35683
rect 33551 35649 33560 35683
rect 33508 35640 33560 35649
rect 31484 35572 31536 35624
rect 29644 35436 29696 35488
rect 29920 35436 29972 35488
rect 30104 35436 30156 35488
rect 31024 35436 31076 35488
rect 32772 35436 32824 35488
rect 33324 35479 33376 35488
rect 33324 35445 33333 35479
rect 33333 35445 33367 35479
rect 33367 35445 33376 35479
rect 33324 35436 33376 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 9772 35232 9824 35284
rect 10968 35232 11020 35284
rect 18880 35232 18932 35284
rect 23480 35232 23532 35284
rect 23940 35232 23992 35284
rect 25412 35232 25464 35284
rect 26516 35232 26568 35284
rect 28172 35275 28224 35284
rect 28172 35241 28181 35275
rect 28181 35241 28215 35275
rect 28215 35241 28224 35275
rect 28172 35232 28224 35241
rect 28356 35232 28408 35284
rect 29920 35232 29972 35284
rect 32772 35232 32824 35284
rect 9864 35164 9916 35216
rect 7196 35096 7248 35148
rect 10784 35164 10836 35216
rect 8208 35028 8260 35080
rect 8300 35028 8352 35080
rect 15108 35096 15160 35148
rect 18788 35096 18840 35148
rect 20996 35096 21048 35148
rect 22560 35096 22612 35148
rect 23664 35139 23716 35148
rect 23664 35105 23673 35139
rect 23673 35105 23707 35139
rect 23707 35105 23716 35139
rect 23664 35096 23716 35105
rect 17316 35071 17368 35080
rect 17316 35037 17325 35071
rect 17325 35037 17359 35071
rect 17359 35037 17368 35071
rect 17316 35028 17368 35037
rect 20812 35028 20864 35080
rect 7196 35003 7248 35012
rect 7196 34969 7205 35003
rect 7205 34969 7239 35003
rect 7239 34969 7248 35003
rect 7196 34960 7248 34969
rect 16120 34960 16172 35012
rect 18144 34960 18196 35012
rect 23572 34960 23624 35012
rect 24860 35164 24912 35216
rect 26148 35164 26200 35216
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 25504 35071 25556 35080
rect 25504 35037 25513 35071
rect 25513 35037 25547 35071
rect 25547 35037 25556 35071
rect 25504 35028 25556 35037
rect 26332 35071 26384 35080
rect 26332 35037 26341 35071
rect 26341 35037 26375 35071
rect 26375 35037 26384 35071
rect 26332 35028 26384 35037
rect 26608 35096 26660 35148
rect 28080 35207 28132 35216
rect 28080 35173 28089 35207
rect 28089 35173 28123 35207
rect 28123 35173 28132 35207
rect 28080 35164 28132 35173
rect 29552 35164 29604 35216
rect 26700 35071 26752 35080
rect 26700 35037 26709 35071
rect 26709 35037 26743 35071
rect 26743 35037 26752 35071
rect 26700 35028 26752 35037
rect 27344 35028 27396 35080
rect 27620 35028 27672 35080
rect 26792 34960 26844 35012
rect 27896 35028 27948 35080
rect 28080 35028 28132 35080
rect 31024 35096 31076 35148
rect 33324 35096 33376 35148
rect 33416 35096 33468 35148
rect 33692 35096 33744 35148
rect 30380 35071 30432 35080
rect 30380 35037 30389 35071
rect 30389 35037 30423 35071
rect 30423 35037 30432 35071
rect 30380 35028 30432 35037
rect 30840 34960 30892 35012
rect 32496 34960 32548 35012
rect 33416 34960 33468 35012
rect 8668 34935 8720 34944
rect 8668 34901 8677 34935
rect 8677 34901 8711 34935
rect 8711 34901 8720 34935
rect 8668 34892 8720 34901
rect 13084 34892 13136 34944
rect 20720 34892 20772 34944
rect 22284 34892 22336 34944
rect 22928 34892 22980 34944
rect 23848 34892 23900 34944
rect 23940 34935 23992 34944
rect 23940 34901 23949 34935
rect 23949 34901 23983 34935
rect 23983 34901 23992 34935
rect 23940 34892 23992 34901
rect 25228 34892 25280 34944
rect 25596 34892 25648 34944
rect 27804 34892 27856 34944
rect 28816 34935 28868 34944
rect 28816 34901 28825 34935
rect 28825 34901 28859 34935
rect 28859 34901 28868 34935
rect 28816 34892 28868 34901
rect 31668 34892 31720 34944
rect 33324 34892 33376 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 7196 34688 7248 34740
rect 5540 34552 5592 34604
rect 11704 34688 11756 34740
rect 13636 34688 13688 34740
rect 17316 34688 17368 34740
rect 17592 34688 17644 34740
rect 8116 34620 8168 34672
rect 16396 34620 16448 34672
rect 16764 34620 16816 34672
rect 20996 34663 21048 34672
rect 20996 34629 21005 34663
rect 21005 34629 21039 34663
rect 21039 34629 21048 34663
rect 20996 34620 21048 34629
rect 21272 34620 21324 34672
rect 8208 34552 8260 34604
rect 11704 34595 11756 34604
rect 11704 34561 11708 34595
rect 11708 34561 11742 34595
rect 11742 34561 11756 34595
rect 11704 34552 11756 34561
rect 11980 34552 12032 34604
rect 8852 34484 8904 34536
rect 12256 34552 12308 34604
rect 17132 34595 17184 34604
rect 8668 34416 8720 34468
rect 11796 34416 11848 34468
rect 5356 34348 5408 34400
rect 8852 34348 8904 34400
rect 9864 34348 9916 34400
rect 11520 34391 11572 34400
rect 11520 34357 11529 34391
rect 11529 34357 11563 34391
rect 11563 34357 11572 34391
rect 11520 34348 11572 34357
rect 17132 34561 17141 34595
rect 17141 34561 17175 34595
rect 17175 34561 17184 34595
rect 17132 34552 17184 34561
rect 22100 34620 22152 34672
rect 22560 34688 22612 34740
rect 23020 34688 23072 34740
rect 23204 34620 23256 34672
rect 14924 34484 14976 34536
rect 14004 34416 14056 34468
rect 22284 34595 22336 34604
rect 22284 34561 22293 34595
rect 22293 34561 22327 34595
rect 22327 34561 22336 34595
rect 22284 34552 22336 34561
rect 12532 34348 12584 34400
rect 13176 34348 13228 34400
rect 16856 34391 16908 34400
rect 16856 34357 16865 34391
rect 16865 34357 16899 34391
rect 16899 34357 16908 34391
rect 16856 34348 16908 34357
rect 16948 34391 17000 34400
rect 16948 34357 16957 34391
rect 16957 34357 16991 34391
rect 16991 34357 17000 34391
rect 16948 34348 17000 34357
rect 17040 34391 17092 34400
rect 17040 34357 17049 34391
rect 17049 34357 17083 34391
rect 17083 34357 17092 34391
rect 17040 34348 17092 34357
rect 18052 34348 18104 34400
rect 20628 34348 20680 34400
rect 23112 34552 23164 34604
rect 23756 34688 23808 34740
rect 25320 34688 25372 34740
rect 26700 34688 26752 34740
rect 28816 34688 28868 34740
rect 30932 34688 30984 34740
rect 31392 34688 31444 34740
rect 33324 34731 33376 34740
rect 23480 34552 23532 34604
rect 23848 34552 23900 34604
rect 25964 34620 26016 34672
rect 26148 34620 26200 34672
rect 28540 34620 28592 34672
rect 33324 34697 33333 34731
rect 33333 34697 33367 34731
rect 33367 34697 33376 34731
rect 33324 34688 33376 34697
rect 33508 34688 33560 34740
rect 26424 34552 26476 34604
rect 31576 34595 31628 34604
rect 31576 34561 31585 34595
rect 31585 34561 31619 34595
rect 31619 34561 31628 34595
rect 31576 34552 31628 34561
rect 31668 34527 31720 34536
rect 31668 34493 31677 34527
rect 31677 34493 31711 34527
rect 31711 34493 31720 34527
rect 31668 34484 31720 34493
rect 24952 34416 25004 34468
rect 26424 34416 26476 34468
rect 30840 34416 30892 34468
rect 31300 34416 31352 34468
rect 32772 34484 32824 34536
rect 36912 34552 36964 34604
rect 34152 34484 34204 34536
rect 37924 34484 37976 34536
rect 22100 34348 22152 34400
rect 22284 34348 22336 34400
rect 23020 34348 23072 34400
rect 23756 34348 23808 34400
rect 24768 34348 24820 34400
rect 27252 34348 27304 34400
rect 28080 34348 28132 34400
rect 29644 34348 29696 34400
rect 30564 34348 30616 34400
rect 30656 34348 30708 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 14832 34187 14884 34196
rect 14832 34153 14841 34187
rect 14841 34153 14875 34187
rect 14875 34153 14884 34187
rect 14832 34144 14884 34153
rect 16488 34144 16540 34196
rect 16856 34144 16908 34196
rect 16948 34144 17000 34196
rect 17132 34144 17184 34196
rect 17316 34144 17368 34196
rect 17960 34144 18012 34196
rect 14280 34076 14332 34128
rect 14372 34076 14424 34128
rect 14464 34076 14516 34128
rect 5724 34008 5776 34060
rect 6368 33940 6420 33992
rect 6828 33940 6880 33992
rect 7288 33983 7340 33992
rect 7288 33949 7297 33983
rect 7297 33949 7331 33983
rect 7331 33949 7340 33983
rect 7288 33940 7340 33949
rect 9036 34008 9088 34060
rect 5356 33872 5408 33924
rect 12072 34008 12124 34060
rect 13176 34051 13228 34060
rect 13176 34017 13185 34051
rect 13185 34017 13219 34051
rect 13219 34017 13228 34051
rect 13176 34008 13228 34017
rect 15384 34051 15436 34060
rect 15384 34017 15393 34051
rect 15393 34017 15427 34051
rect 15427 34017 15436 34051
rect 15384 34008 15436 34017
rect 16856 34051 16908 34060
rect 16856 34017 16865 34051
rect 16865 34017 16899 34051
rect 16899 34017 16908 34051
rect 16856 34008 16908 34017
rect 17776 34076 17828 34128
rect 20536 34076 20588 34128
rect 9864 33983 9916 33992
rect 9864 33949 9873 33983
rect 9873 33949 9907 33983
rect 9907 33949 9916 33983
rect 9864 33940 9916 33949
rect 11520 33940 11572 33992
rect 11796 33983 11848 33992
rect 11796 33949 11805 33983
rect 11805 33949 11839 33983
rect 11839 33949 11848 33983
rect 11796 33940 11848 33949
rect 6736 33847 6788 33856
rect 6736 33813 6745 33847
rect 6745 33813 6779 33847
rect 6779 33813 6788 33847
rect 9588 33872 9640 33924
rect 13360 33940 13412 33992
rect 14464 33940 14516 33992
rect 16028 33983 16080 33992
rect 16028 33949 16037 33983
rect 16037 33949 16071 33983
rect 16071 33949 16080 33983
rect 16028 33940 16080 33949
rect 16212 33983 16264 33992
rect 16212 33949 16221 33983
rect 16221 33949 16255 33983
rect 16255 33949 16264 33983
rect 16212 33940 16264 33949
rect 16304 33983 16356 33992
rect 16304 33949 16313 33983
rect 16313 33949 16347 33983
rect 16347 33949 16356 33983
rect 16304 33940 16356 33949
rect 16396 33983 16448 33992
rect 16396 33949 16405 33983
rect 16405 33949 16439 33983
rect 16439 33949 16448 33983
rect 16396 33940 16448 33949
rect 17132 33940 17184 33992
rect 17316 33940 17368 33992
rect 17684 33983 17736 33992
rect 17684 33949 17693 33983
rect 17693 33949 17727 33983
rect 17727 33949 17736 33983
rect 17684 33940 17736 33949
rect 6736 33804 6788 33813
rect 7196 33847 7248 33856
rect 7196 33813 7205 33847
rect 7205 33813 7239 33847
rect 7239 33813 7248 33847
rect 7196 33804 7248 33813
rect 8668 33847 8720 33856
rect 8668 33813 8677 33847
rect 8677 33813 8711 33847
rect 8711 33813 8720 33847
rect 8668 33804 8720 33813
rect 8944 33847 8996 33856
rect 8944 33813 8953 33847
rect 8953 33813 8987 33847
rect 8987 33813 8996 33847
rect 8944 33804 8996 33813
rect 9404 33804 9456 33856
rect 11888 33804 11940 33856
rect 13268 33804 13320 33856
rect 13728 33804 13780 33856
rect 14556 33804 14608 33856
rect 14648 33804 14700 33856
rect 15660 33847 15712 33856
rect 15660 33813 15669 33847
rect 15669 33813 15703 33847
rect 15703 33813 15712 33847
rect 15660 33804 15712 33813
rect 16028 33804 16080 33856
rect 16396 33804 16448 33856
rect 17960 33915 18012 33924
rect 17960 33881 17969 33915
rect 17969 33881 18003 33915
rect 18003 33881 18012 33915
rect 17960 33872 18012 33881
rect 18052 33915 18104 33924
rect 18052 33881 18061 33915
rect 18061 33881 18095 33915
rect 18095 33881 18104 33915
rect 18052 33872 18104 33881
rect 16948 33804 17000 33856
rect 17137 33847 17189 33856
rect 17137 33813 17141 33847
rect 17141 33813 17175 33847
rect 17175 33813 17189 33847
rect 17137 33804 17189 33813
rect 17316 33804 17368 33856
rect 18420 33983 18472 33992
rect 18420 33949 18429 33983
rect 18429 33949 18463 33983
rect 18463 33949 18472 33983
rect 18420 33940 18472 33949
rect 18236 33872 18288 33924
rect 18604 33915 18656 33924
rect 18604 33881 18613 33915
rect 18613 33881 18647 33915
rect 18647 33881 18656 33915
rect 18604 33872 18656 33881
rect 18788 33983 18840 33992
rect 18788 33949 18797 33983
rect 18797 33949 18831 33983
rect 18831 33949 18840 33983
rect 18788 33940 18840 33949
rect 19248 33983 19300 33992
rect 19248 33949 19257 33983
rect 19257 33949 19291 33983
rect 19291 33949 19300 33983
rect 19248 33940 19300 33949
rect 19064 33872 19116 33924
rect 18328 33847 18380 33856
rect 18328 33813 18337 33847
rect 18337 33813 18371 33847
rect 18371 33813 18380 33847
rect 18328 33804 18380 33813
rect 20260 33983 20312 33992
rect 20260 33949 20269 33983
rect 20269 33949 20303 33983
rect 20303 33949 20312 33983
rect 20260 33940 20312 33949
rect 20536 33940 20588 33992
rect 20628 33940 20680 33992
rect 21732 33940 21784 33992
rect 21916 33983 21968 33992
rect 21916 33949 21925 33983
rect 21925 33949 21959 33983
rect 21959 33949 21968 33983
rect 21916 33940 21968 33949
rect 22100 33983 22152 33992
rect 22100 33949 22109 33983
rect 22109 33949 22143 33983
rect 22143 33949 22152 33983
rect 22100 33940 22152 33949
rect 22284 33940 22336 33992
rect 22468 33940 22520 33992
rect 20352 33804 20404 33856
rect 21732 33804 21784 33856
rect 22468 33804 22520 33856
rect 22560 33804 22612 33856
rect 23204 33983 23256 33992
rect 23204 33949 23213 33983
rect 23213 33949 23247 33983
rect 23247 33949 23256 33983
rect 23204 33940 23256 33949
rect 23480 33983 23532 33992
rect 23480 33949 23489 33983
rect 23489 33949 23523 33983
rect 23523 33949 23532 33983
rect 23480 33940 23532 33949
rect 23572 33983 23624 33992
rect 23572 33949 23581 33983
rect 23581 33949 23615 33983
rect 23615 33949 23624 33983
rect 23572 33940 23624 33949
rect 24216 33940 24268 33992
rect 24768 33940 24820 33992
rect 25412 33940 25464 33992
rect 24032 33872 24084 33924
rect 23020 33804 23072 33856
rect 23112 33847 23164 33856
rect 23112 33813 23121 33847
rect 23121 33813 23155 33847
rect 23155 33813 23164 33847
rect 23112 33804 23164 33813
rect 23848 33847 23900 33856
rect 23848 33813 23857 33847
rect 23857 33813 23891 33847
rect 23891 33813 23900 33847
rect 23848 33804 23900 33813
rect 24492 33804 24544 33856
rect 25412 33847 25464 33856
rect 25412 33813 25421 33847
rect 25421 33813 25455 33847
rect 25455 33813 25464 33847
rect 25412 33804 25464 33813
rect 28080 34187 28132 34196
rect 28080 34153 28089 34187
rect 28089 34153 28123 34187
rect 28123 34153 28132 34187
rect 28080 34144 28132 34153
rect 30840 34144 30892 34196
rect 25964 33983 26016 33992
rect 25964 33949 25973 33983
rect 25973 33949 26007 33983
rect 26007 33949 26016 33983
rect 25964 33940 26016 33949
rect 26148 33940 26200 33992
rect 28448 34119 28500 34128
rect 28448 34085 28457 34119
rect 28457 34085 28491 34119
rect 28491 34085 28500 34119
rect 28448 34076 28500 34085
rect 26424 33915 26476 33924
rect 26424 33881 26433 33915
rect 26433 33881 26467 33915
rect 26467 33881 26476 33915
rect 26424 33872 26476 33881
rect 26976 33940 27028 33992
rect 28448 33940 28500 33992
rect 28632 33940 28684 33992
rect 27160 33847 27212 33856
rect 27160 33813 27169 33847
rect 27169 33813 27203 33847
rect 27203 33813 27212 33847
rect 27160 33804 27212 33813
rect 28172 33804 28224 33856
rect 28816 33847 28868 33856
rect 28816 33813 28825 33847
rect 28825 33813 28859 33847
rect 28859 33813 28868 33847
rect 28816 33804 28868 33813
rect 29644 33804 29696 33856
rect 29920 34076 29972 34128
rect 29828 33940 29880 33992
rect 30472 33983 30524 33992
rect 30472 33949 30481 33983
rect 30481 33949 30515 33983
rect 30515 33949 30524 33983
rect 30472 33940 30524 33949
rect 30564 33983 30616 33992
rect 30564 33949 30574 33983
rect 30574 33949 30608 33983
rect 30608 33949 30616 33983
rect 30564 33940 30616 33949
rect 30840 33983 30892 33992
rect 30840 33949 30849 33983
rect 30849 33949 30883 33983
rect 30883 33949 30892 33983
rect 30840 33940 30892 33949
rect 31484 33983 31536 33992
rect 31484 33949 31493 33983
rect 31493 33949 31527 33983
rect 31527 33949 31536 33983
rect 31484 33940 31536 33949
rect 33876 33983 33928 33992
rect 33876 33949 33885 33983
rect 33885 33949 33919 33983
rect 33919 33949 33928 33983
rect 33876 33940 33928 33949
rect 34336 33983 34388 33992
rect 34336 33949 34345 33983
rect 34345 33949 34379 33983
rect 34379 33949 34388 33983
rect 34336 33940 34388 33949
rect 31668 33804 31720 33856
rect 32220 33804 32272 33856
rect 33324 33804 33376 33856
rect 36268 33872 36320 33924
rect 35992 33804 36044 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 5540 33600 5592 33652
rect 6736 33600 6788 33652
rect 7196 33600 7248 33652
rect 8668 33600 8720 33652
rect 8300 33464 8352 33516
rect 9404 33600 9456 33652
rect 13360 33600 13412 33652
rect 13912 33600 13964 33652
rect 14648 33600 14700 33652
rect 16672 33600 16724 33652
rect 17316 33600 17368 33652
rect 17684 33600 17736 33652
rect 19340 33600 19392 33652
rect 11796 33532 11848 33584
rect 10324 33464 10376 33516
rect 5908 33439 5960 33448
rect 5908 33405 5917 33439
rect 5917 33405 5951 33439
rect 5951 33405 5960 33439
rect 5908 33396 5960 33405
rect 7288 33439 7340 33448
rect 7288 33405 7297 33439
rect 7297 33405 7331 33439
rect 7331 33405 7340 33439
rect 7288 33396 7340 33405
rect 9588 33396 9640 33448
rect 16488 33532 16540 33584
rect 13268 33464 13320 33516
rect 13544 33464 13596 33516
rect 14004 33439 14056 33448
rect 14004 33405 14013 33439
rect 14013 33405 14047 33439
rect 14047 33405 14056 33439
rect 14004 33396 14056 33405
rect 15752 33328 15804 33380
rect 7472 33260 7524 33312
rect 10600 33260 10652 33312
rect 11796 33260 11848 33312
rect 16212 33260 16264 33312
rect 17776 33464 17828 33516
rect 19708 33507 19760 33516
rect 19708 33473 19742 33507
rect 19742 33473 19760 33507
rect 19708 33464 19760 33473
rect 20260 33600 20312 33652
rect 21088 33643 21140 33652
rect 21088 33609 21097 33643
rect 21097 33609 21131 33643
rect 21131 33609 21140 33643
rect 21088 33600 21140 33609
rect 21272 33643 21324 33652
rect 21272 33609 21281 33643
rect 21281 33609 21315 33643
rect 21315 33609 21324 33643
rect 21272 33600 21324 33609
rect 21916 33600 21968 33652
rect 22468 33600 22520 33652
rect 22652 33600 22704 33652
rect 22836 33600 22888 33652
rect 23020 33600 23072 33652
rect 27160 33600 27212 33652
rect 27344 33600 27396 33652
rect 20352 33507 20404 33516
rect 20352 33473 20361 33507
rect 20361 33473 20395 33507
rect 20395 33473 20404 33507
rect 20352 33464 20404 33473
rect 20628 33507 20680 33516
rect 20628 33473 20637 33507
rect 20637 33473 20671 33507
rect 20671 33473 20680 33507
rect 20628 33464 20680 33473
rect 19064 33439 19116 33448
rect 19064 33405 19073 33439
rect 19073 33405 19107 33439
rect 19107 33405 19116 33439
rect 19064 33396 19116 33405
rect 19616 33396 19668 33448
rect 21456 33575 21508 33584
rect 21456 33541 21465 33575
rect 21465 33541 21499 33575
rect 21499 33541 21508 33575
rect 21456 33532 21508 33541
rect 23296 33532 23348 33584
rect 20812 33396 20864 33448
rect 21824 33507 21876 33516
rect 21824 33473 21833 33507
rect 21833 33473 21867 33507
rect 21867 33473 21876 33507
rect 21824 33464 21876 33473
rect 23756 33507 23808 33516
rect 23756 33473 23765 33507
rect 23765 33473 23799 33507
rect 23799 33473 23808 33507
rect 23756 33464 23808 33473
rect 23848 33507 23900 33516
rect 23848 33473 23857 33507
rect 23857 33473 23891 33507
rect 23891 33473 23900 33507
rect 23848 33464 23900 33473
rect 25320 33532 25372 33584
rect 23480 33439 23532 33448
rect 23480 33405 23489 33439
rect 23489 33405 23523 33439
rect 23523 33405 23532 33439
rect 23480 33396 23532 33405
rect 23940 33396 23992 33448
rect 25412 33396 25464 33448
rect 17592 33328 17644 33380
rect 18144 33328 18196 33380
rect 19892 33328 19944 33380
rect 19984 33328 20036 33380
rect 18420 33260 18472 33312
rect 19432 33260 19484 33312
rect 20536 33260 20588 33312
rect 21456 33260 21508 33312
rect 22100 33260 22152 33312
rect 23848 33260 23900 33312
rect 24032 33303 24084 33312
rect 24032 33269 24041 33303
rect 24041 33269 24075 33303
rect 24075 33269 24084 33303
rect 24032 33260 24084 33269
rect 25412 33303 25464 33312
rect 25412 33269 25421 33303
rect 25421 33269 25455 33303
rect 25455 33269 25464 33303
rect 25412 33260 25464 33269
rect 26608 33507 26660 33516
rect 26608 33473 26617 33507
rect 26617 33473 26651 33507
rect 26651 33473 26660 33507
rect 26608 33464 26660 33473
rect 28540 33532 28592 33584
rect 28816 33532 28868 33584
rect 31576 33532 31628 33584
rect 33140 33600 33192 33652
rect 33876 33600 33928 33652
rect 34152 33643 34204 33652
rect 34152 33609 34161 33643
rect 34161 33609 34195 33643
rect 34195 33609 34204 33643
rect 34152 33600 34204 33609
rect 29184 33464 29236 33516
rect 33324 33464 33376 33516
rect 27804 33396 27856 33448
rect 34060 33439 34112 33448
rect 34060 33405 34069 33439
rect 34069 33405 34103 33439
rect 34103 33405 34112 33439
rect 34060 33396 34112 33405
rect 34244 33507 34296 33516
rect 34244 33473 34253 33507
rect 34253 33473 34287 33507
rect 34287 33473 34296 33507
rect 34244 33464 34296 33473
rect 36912 33643 36964 33652
rect 36912 33609 36921 33643
rect 36921 33609 36955 33643
rect 36955 33609 36964 33643
rect 36912 33600 36964 33609
rect 36268 33464 36320 33516
rect 36728 33507 36780 33516
rect 36728 33473 36737 33507
rect 36737 33473 36771 33507
rect 36771 33473 36780 33507
rect 36728 33464 36780 33473
rect 33232 33260 33284 33312
rect 34244 33260 34296 33312
rect 34796 33260 34848 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 3976 32852 4028 32904
rect 7196 33056 7248 33108
rect 7288 33056 7340 33108
rect 8944 33056 8996 33108
rect 6368 32988 6420 33040
rect 5908 32852 5960 32904
rect 6552 32852 6604 32904
rect 4896 32784 4948 32836
rect 6828 32963 6880 32972
rect 6828 32929 6837 32963
rect 6837 32929 6871 32963
rect 6871 32929 6880 32963
rect 6828 32920 6880 32929
rect 7840 32895 7892 32904
rect 7840 32861 7849 32895
rect 7849 32861 7883 32895
rect 7883 32861 7892 32895
rect 7840 32852 7892 32861
rect 9772 33056 9824 33108
rect 9864 33056 9916 33108
rect 17316 33056 17368 33108
rect 18328 33056 18380 33108
rect 8208 32895 8260 32904
rect 8208 32861 8217 32895
rect 8217 32861 8251 32895
rect 8251 32861 8260 32895
rect 8208 32852 8260 32861
rect 8116 32784 8168 32836
rect 6276 32759 6328 32768
rect 6276 32725 6285 32759
rect 6285 32725 6319 32759
rect 6319 32725 6328 32759
rect 6276 32716 6328 32725
rect 7380 32716 7432 32768
rect 8576 32852 8628 32904
rect 12624 32988 12676 33040
rect 20536 33056 20588 33108
rect 24492 33056 24544 33108
rect 26608 33099 26660 33108
rect 26608 33065 26617 33099
rect 26617 33065 26651 33099
rect 26651 33065 26660 33099
rect 26608 33056 26660 33065
rect 29552 33056 29604 33108
rect 30472 33056 30524 33108
rect 30656 33056 30708 33108
rect 31300 33056 31352 33108
rect 33324 33056 33376 33108
rect 34796 33056 34848 33108
rect 10600 32852 10652 32904
rect 11520 32852 11572 32904
rect 11796 32852 11848 32904
rect 18880 32920 18932 32972
rect 19616 32963 19668 32972
rect 19616 32929 19629 32963
rect 19629 32929 19663 32963
rect 19663 32929 19668 32963
rect 19616 32920 19668 32929
rect 20168 32988 20220 33040
rect 11980 32827 12032 32836
rect 11980 32793 11989 32827
rect 11989 32793 12023 32827
rect 12023 32793 12032 32827
rect 11980 32784 12032 32793
rect 12072 32827 12124 32836
rect 12072 32793 12081 32827
rect 12081 32793 12115 32827
rect 12115 32793 12124 32827
rect 12072 32784 12124 32793
rect 8852 32716 8904 32768
rect 9772 32716 9824 32768
rect 10508 32716 10560 32768
rect 11796 32716 11848 32768
rect 15752 32852 15804 32904
rect 15844 32852 15896 32904
rect 16212 32895 16264 32904
rect 16212 32861 16221 32895
rect 16221 32861 16255 32895
rect 16255 32861 16264 32895
rect 16212 32852 16264 32861
rect 16396 32852 16448 32904
rect 17224 32852 17276 32904
rect 18696 32895 18748 32904
rect 18696 32861 18705 32895
rect 18705 32861 18739 32895
rect 18739 32861 18748 32895
rect 18696 32852 18748 32861
rect 18236 32784 18288 32836
rect 12348 32759 12400 32768
rect 12348 32725 12357 32759
rect 12357 32725 12391 32759
rect 12391 32725 12400 32759
rect 12348 32716 12400 32725
rect 16672 32716 16724 32768
rect 19064 32784 19116 32836
rect 19708 32852 19760 32904
rect 20260 32852 20312 32904
rect 22008 32988 22060 33040
rect 26148 32988 26200 33040
rect 20536 32895 20588 32904
rect 20536 32861 20545 32895
rect 20545 32861 20579 32895
rect 20579 32861 20588 32895
rect 20536 32852 20588 32861
rect 20904 32852 20956 32904
rect 21456 32895 21508 32904
rect 21456 32861 21465 32895
rect 21465 32861 21499 32895
rect 21499 32861 21508 32895
rect 21456 32852 21508 32861
rect 19984 32784 20036 32836
rect 26884 32920 26936 32972
rect 21916 32852 21968 32904
rect 22192 32852 22244 32904
rect 22836 32852 22888 32904
rect 27804 32920 27856 32972
rect 28540 32920 28592 32972
rect 20720 32759 20772 32768
rect 20720 32725 20729 32759
rect 20729 32725 20763 32759
rect 20763 32725 20772 32759
rect 20720 32716 20772 32725
rect 21548 32716 21600 32768
rect 23940 32716 23992 32768
rect 26332 32716 26384 32768
rect 26608 32716 26660 32768
rect 27528 32895 27580 32904
rect 27528 32861 27537 32895
rect 27537 32861 27571 32895
rect 27571 32861 27580 32895
rect 27528 32852 27580 32861
rect 28816 32852 28868 32904
rect 30288 32852 30340 32904
rect 30932 32895 30984 32904
rect 30932 32861 30941 32895
rect 30941 32861 30975 32895
rect 30975 32861 30984 32895
rect 30932 32852 30984 32861
rect 31208 32895 31260 32904
rect 31208 32861 31217 32895
rect 31217 32861 31251 32895
rect 31251 32861 31260 32895
rect 31208 32852 31260 32861
rect 32496 32852 32548 32904
rect 32956 32852 33008 32904
rect 34336 32895 34388 32904
rect 34336 32861 34345 32895
rect 34345 32861 34379 32895
rect 34379 32861 34388 32895
rect 34336 32852 34388 32861
rect 35992 32852 36044 32904
rect 28080 32784 28132 32836
rect 29092 32784 29144 32836
rect 27252 32716 27304 32768
rect 27620 32716 27672 32768
rect 28724 32716 28776 32768
rect 30196 32759 30248 32768
rect 30196 32725 30205 32759
rect 30205 32725 30239 32759
rect 30239 32725 30248 32759
rect 30196 32716 30248 32725
rect 32128 32716 32180 32768
rect 35624 32716 35676 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4896 32512 4948 32564
rect 6276 32512 6328 32564
rect 8116 32512 8168 32564
rect 12348 32512 12400 32564
rect 17684 32555 17736 32564
rect 17684 32521 17693 32555
rect 17693 32521 17727 32555
rect 17727 32521 17736 32555
rect 17684 32512 17736 32521
rect 5724 32308 5776 32360
rect 8300 32308 8352 32360
rect 11888 32419 11940 32428
rect 11888 32385 11897 32419
rect 11897 32385 11931 32419
rect 11931 32385 11940 32419
rect 11888 32376 11940 32385
rect 16396 32444 16448 32496
rect 17040 32444 17092 32496
rect 17500 32487 17552 32496
rect 17500 32453 17509 32487
rect 17509 32453 17543 32487
rect 17543 32453 17552 32487
rect 17500 32444 17552 32453
rect 13544 32376 13596 32428
rect 20260 32444 20312 32496
rect 21640 32444 21692 32496
rect 16120 32308 16172 32360
rect 12256 32240 12308 32292
rect 13636 32240 13688 32292
rect 18420 32419 18472 32428
rect 18420 32385 18429 32419
rect 18429 32385 18463 32419
rect 18463 32385 18472 32419
rect 18420 32376 18472 32385
rect 18604 32419 18656 32428
rect 18604 32385 18613 32419
rect 18613 32385 18647 32419
rect 18647 32385 18656 32419
rect 18604 32376 18656 32385
rect 18696 32419 18748 32428
rect 18696 32385 18705 32419
rect 18705 32385 18739 32419
rect 18739 32385 18748 32419
rect 18696 32376 18748 32385
rect 18972 32419 19024 32428
rect 18972 32385 18981 32419
rect 18981 32385 19015 32419
rect 19015 32385 19024 32419
rect 18972 32376 19024 32385
rect 19064 32376 19116 32428
rect 17592 32240 17644 32292
rect 21272 32419 21324 32428
rect 21272 32385 21281 32419
rect 21281 32385 21315 32419
rect 21315 32385 21324 32419
rect 21272 32376 21324 32385
rect 21364 32376 21416 32428
rect 22284 32376 22336 32428
rect 23388 32512 23440 32564
rect 23848 32512 23900 32564
rect 22836 32444 22888 32496
rect 23296 32444 23348 32496
rect 23388 32419 23440 32428
rect 23388 32385 23397 32419
rect 23397 32385 23431 32419
rect 23431 32385 23440 32419
rect 23388 32376 23440 32385
rect 23940 32487 23992 32496
rect 23940 32453 23949 32487
rect 23949 32453 23983 32487
rect 23983 32453 23992 32487
rect 23940 32444 23992 32453
rect 27528 32512 27580 32564
rect 28080 32512 28132 32564
rect 31208 32512 31260 32564
rect 36728 32512 36780 32564
rect 27712 32444 27764 32496
rect 23112 32308 23164 32360
rect 24124 32419 24176 32428
rect 24124 32385 24133 32419
rect 24133 32385 24167 32419
rect 24167 32385 24176 32419
rect 24124 32376 24176 32385
rect 25964 32376 26016 32428
rect 24768 32308 24820 32360
rect 25780 32308 25832 32360
rect 11612 32172 11664 32224
rect 15660 32172 15712 32224
rect 16764 32172 16816 32224
rect 17132 32172 17184 32224
rect 19432 32172 19484 32224
rect 19984 32215 20036 32224
rect 19984 32181 19993 32215
rect 19993 32181 20027 32215
rect 20027 32181 20036 32215
rect 19984 32172 20036 32181
rect 22192 32215 22244 32224
rect 22192 32181 22201 32215
rect 22201 32181 22235 32215
rect 22235 32181 22244 32215
rect 22192 32172 22244 32181
rect 22836 32215 22888 32224
rect 22836 32181 22845 32215
rect 22845 32181 22879 32215
rect 22879 32181 22888 32215
rect 22836 32172 22888 32181
rect 25320 32172 25372 32224
rect 27988 32308 28040 32360
rect 28356 32308 28408 32360
rect 28448 32351 28500 32360
rect 28448 32317 28457 32351
rect 28457 32317 28491 32351
rect 28491 32317 28500 32351
rect 28448 32308 28500 32317
rect 26700 32240 26752 32292
rect 28724 32376 28776 32428
rect 30656 32351 30708 32360
rect 30656 32317 30665 32351
rect 30665 32317 30699 32351
rect 30699 32317 30708 32351
rect 30656 32308 30708 32317
rect 30840 32419 30892 32428
rect 30840 32385 30849 32419
rect 30849 32385 30883 32419
rect 30883 32385 30892 32419
rect 30840 32376 30892 32385
rect 32588 32444 32640 32496
rect 34612 32444 34664 32496
rect 32128 32376 32180 32428
rect 32220 32376 32272 32428
rect 33140 32419 33192 32428
rect 33140 32385 33149 32419
rect 33149 32385 33183 32419
rect 33183 32385 33192 32419
rect 33140 32376 33192 32385
rect 33232 32376 33284 32428
rect 35624 32419 35676 32428
rect 35624 32385 35633 32419
rect 35633 32385 35667 32419
rect 35667 32385 35676 32419
rect 35624 32376 35676 32385
rect 32312 32308 32364 32360
rect 30932 32240 30984 32292
rect 32864 32283 32916 32292
rect 32864 32249 32873 32283
rect 32873 32249 32907 32283
rect 32907 32249 32916 32283
rect 32864 32240 32916 32249
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 7840 31968 7892 32020
rect 8576 31968 8628 32020
rect 13544 31968 13596 32020
rect 17592 31968 17644 32020
rect 18144 31968 18196 32020
rect 18972 31968 19024 32020
rect 19064 32011 19116 32020
rect 19064 31977 19073 32011
rect 19073 31977 19107 32011
rect 19107 31977 19116 32011
rect 19064 31968 19116 31977
rect 22008 31968 22060 32020
rect 22560 31968 22612 32020
rect 5724 31832 5776 31884
rect 11612 31900 11664 31952
rect 3976 31807 4028 31816
rect 3976 31773 3985 31807
rect 3985 31773 4019 31807
rect 4019 31773 4028 31807
rect 3976 31764 4028 31773
rect 6552 31764 6604 31816
rect 7380 31764 7432 31816
rect 7656 31807 7708 31816
rect 7656 31773 7665 31807
rect 7665 31773 7699 31807
rect 7699 31773 7708 31807
rect 7656 31764 7708 31773
rect 9036 31832 9088 31884
rect 8116 31807 8168 31816
rect 8116 31773 8125 31807
rect 8125 31773 8159 31807
rect 8159 31773 8168 31807
rect 8116 31764 8168 31773
rect 8484 31807 8536 31816
rect 8484 31773 8493 31807
rect 8493 31773 8527 31807
rect 8527 31773 8536 31807
rect 8484 31764 8536 31773
rect 8852 31764 8904 31816
rect 17960 31832 18012 31884
rect 18328 31832 18380 31884
rect 20352 31900 20404 31952
rect 21824 31900 21876 31952
rect 14464 31764 14516 31816
rect 15476 31764 15528 31816
rect 16396 31764 16448 31816
rect 20628 31832 20680 31884
rect 22744 31900 22796 31952
rect 23020 31900 23072 31952
rect 23112 31900 23164 31952
rect 23388 31900 23440 31952
rect 9772 31739 9824 31748
rect 9772 31705 9781 31739
rect 9781 31705 9815 31739
rect 9815 31705 9824 31739
rect 9772 31696 9824 31705
rect 10324 31696 10376 31748
rect 12900 31696 12952 31748
rect 13268 31739 13320 31748
rect 13268 31705 13277 31739
rect 13277 31705 13311 31739
rect 13311 31705 13320 31739
rect 13268 31696 13320 31705
rect 7840 31628 7892 31680
rect 8300 31671 8352 31680
rect 8300 31637 8309 31671
rect 8309 31637 8343 31671
rect 8343 31637 8352 31671
rect 8300 31628 8352 31637
rect 11612 31628 11664 31680
rect 13360 31671 13412 31680
rect 13360 31637 13369 31671
rect 13369 31637 13403 31671
rect 13403 31637 13412 31671
rect 13360 31628 13412 31637
rect 13912 31696 13964 31748
rect 21272 31807 21324 31816
rect 21272 31773 21281 31807
rect 21281 31773 21315 31807
rect 21315 31773 21324 31807
rect 21272 31764 21324 31773
rect 21916 31807 21968 31816
rect 21916 31773 21925 31807
rect 21925 31773 21959 31807
rect 21959 31773 21968 31807
rect 21916 31764 21968 31773
rect 22008 31807 22060 31816
rect 22008 31773 22018 31807
rect 22018 31773 22052 31807
rect 22052 31773 22060 31807
rect 22008 31764 22060 31773
rect 22100 31764 22152 31816
rect 22376 31807 22428 31816
rect 22376 31773 22390 31807
rect 22390 31773 22424 31807
rect 22424 31773 22428 31807
rect 22376 31764 22428 31773
rect 17224 31696 17276 31748
rect 20536 31696 20588 31748
rect 23112 31807 23164 31816
rect 23112 31773 23126 31807
rect 23126 31773 23160 31807
rect 23160 31773 23164 31807
rect 23112 31764 23164 31773
rect 23296 31764 23348 31816
rect 24124 31832 24176 31884
rect 23572 31764 23624 31816
rect 23664 31807 23716 31816
rect 23664 31773 23673 31807
rect 23673 31773 23707 31807
rect 23707 31773 23716 31807
rect 23664 31764 23716 31773
rect 23940 31764 23992 31816
rect 24216 31764 24268 31816
rect 24308 31764 24360 31816
rect 25136 31968 25188 32020
rect 24584 31832 24636 31884
rect 25504 31900 25556 31952
rect 26976 31900 27028 31952
rect 28724 31900 28776 31952
rect 22928 31739 22980 31748
rect 22928 31705 22937 31739
rect 22937 31705 22971 31739
rect 22971 31705 22980 31739
rect 22928 31696 22980 31705
rect 23756 31739 23808 31748
rect 23756 31705 23765 31739
rect 23765 31705 23799 31739
rect 23799 31705 23808 31739
rect 23756 31696 23808 31705
rect 25044 31764 25096 31816
rect 25136 31807 25188 31816
rect 25136 31773 25145 31807
rect 25145 31773 25179 31807
rect 25179 31773 25188 31807
rect 25136 31764 25188 31773
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 26056 31764 26108 31816
rect 26700 31764 26752 31816
rect 29092 31832 29144 31884
rect 27896 31764 27948 31816
rect 28264 31807 28316 31816
rect 28264 31773 28273 31807
rect 28273 31773 28307 31807
rect 28307 31773 28316 31807
rect 28264 31764 28316 31773
rect 29276 31764 29328 31816
rect 29552 31807 29604 31816
rect 29552 31773 29561 31807
rect 29561 31773 29595 31807
rect 29595 31773 29604 31807
rect 29552 31764 29604 31773
rect 18144 31628 18196 31680
rect 18696 31671 18748 31680
rect 18696 31637 18705 31671
rect 18705 31637 18739 31671
rect 18739 31637 18748 31671
rect 18696 31628 18748 31637
rect 20168 31628 20220 31680
rect 22560 31671 22612 31680
rect 22560 31637 22569 31671
rect 22569 31637 22603 31671
rect 22603 31637 22612 31671
rect 22560 31628 22612 31637
rect 22652 31628 22704 31680
rect 22744 31628 22796 31680
rect 23388 31628 23440 31680
rect 24768 31628 24820 31680
rect 24952 31628 25004 31680
rect 27344 31696 27396 31748
rect 25596 31671 25648 31680
rect 25596 31637 25605 31671
rect 25605 31637 25639 31671
rect 25639 31637 25648 31671
rect 25596 31628 25648 31637
rect 25780 31628 25832 31680
rect 26148 31628 26200 31680
rect 27712 31628 27764 31680
rect 27988 31628 28040 31680
rect 29552 31628 29604 31680
rect 29828 31807 29880 31816
rect 29828 31773 29837 31807
rect 29837 31773 29871 31807
rect 29871 31773 29880 31807
rect 29828 31764 29880 31773
rect 30288 31832 30340 31884
rect 30012 31807 30064 31816
rect 30012 31773 30026 31807
rect 30026 31773 30060 31807
rect 30060 31773 30064 31807
rect 30012 31764 30064 31773
rect 31484 31807 31536 31816
rect 31484 31773 31493 31807
rect 31493 31773 31527 31807
rect 31527 31773 31536 31807
rect 31484 31764 31536 31773
rect 32128 31968 32180 32020
rect 34612 31764 34664 31816
rect 35440 31807 35492 31816
rect 35440 31773 35449 31807
rect 35449 31773 35483 31807
rect 35483 31773 35492 31807
rect 35440 31764 35492 31773
rect 34520 31696 34572 31748
rect 30380 31671 30432 31680
rect 30380 31637 30389 31671
rect 30389 31637 30423 31671
rect 30423 31637 30432 31671
rect 30380 31628 30432 31637
rect 30748 31628 30800 31680
rect 32036 31628 32088 31680
rect 34796 31671 34848 31680
rect 34796 31637 34805 31671
rect 34805 31637 34839 31671
rect 34839 31637 34848 31671
rect 34796 31628 34848 31637
rect 35256 31671 35308 31680
rect 35256 31637 35265 31671
rect 35265 31637 35299 31671
rect 35299 31637 35308 31671
rect 35256 31628 35308 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 8300 31424 8352 31476
rect 8944 31424 8996 31476
rect 9496 31424 9548 31476
rect 9772 31424 9824 31476
rect 8392 31356 8444 31408
rect 10508 31424 10560 31476
rect 10968 31424 11020 31476
rect 13452 31467 13504 31476
rect 13452 31433 13461 31467
rect 13461 31433 13495 31467
rect 13495 31433 13504 31467
rect 13452 31424 13504 31433
rect 11980 31356 12032 31408
rect 12532 31356 12584 31408
rect 16672 31424 16724 31476
rect 18604 31424 18656 31476
rect 18696 31467 18748 31476
rect 18696 31433 18705 31467
rect 18705 31433 18739 31467
rect 18739 31433 18748 31467
rect 18696 31424 18748 31433
rect 21180 31424 21232 31476
rect 21364 31424 21416 31476
rect 21456 31424 21508 31476
rect 22192 31467 22244 31476
rect 22192 31433 22201 31467
rect 22201 31433 22235 31467
rect 22235 31433 22244 31467
rect 22192 31424 22244 31433
rect 23296 31424 23348 31476
rect 27620 31424 27672 31476
rect 30380 31424 30432 31476
rect 34796 31424 34848 31476
rect 11612 31288 11664 31340
rect 7840 31263 7892 31272
rect 7840 31229 7849 31263
rect 7849 31229 7883 31263
rect 7883 31229 7892 31263
rect 7840 31220 7892 31229
rect 10232 31220 10284 31272
rect 10968 31220 11020 31272
rect 11888 31331 11940 31340
rect 11888 31297 11897 31331
rect 11897 31297 11931 31331
rect 11931 31297 11940 31331
rect 11888 31288 11940 31297
rect 12348 31288 12400 31340
rect 15844 31356 15896 31408
rect 16120 31399 16172 31408
rect 16120 31365 16129 31399
rect 16129 31365 16163 31399
rect 16163 31365 16172 31399
rect 16120 31356 16172 31365
rect 16396 31356 16448 31408
rect 15476 31331 15528 31340
rect 15476 31297 15485 31331
rect 15485 31297 15519 31331
rect 15519 31297 15528 31331
rect 15476 31288 15528 31297
rect 15752 31288 15804 31340
rect 16028 31288 16080 31340
rect 16212 31331 16264 31340
rect 16212 31297 16221 31331
rect 16221 31297 16255 31331
rect 16255 31297 16264 31331
rect 16212 31288 16264 31297
rect 9588 31195 9640 31204
rect 9588 31161 9597 31195
rect 9597 31161 9631 31195
rect 9631 31161 9640 31195
rect 12900 31220 12952 31272
rect 9588 31152 9640 31161
rect 16212 31152 16264 31204
rect 13544 31084 13596 31136
rect 14648 31084 14700 31136
rect 16488 31127 16540 31136
rect 16488 31093 16497 31127
rect 16497 31093 16531 31127
rect 16531 31093 16540 31127
rect 16488 31084 16540 31093
rect 16672 31152 16724 31204
rect 17316 31288 17368 31340
rect 17224 31152 17276 31204
rect 17868 31356 17920 31408
rect 19984 31356 20036 31408
rect 25504 31356 25556 31408
rect 27988 31399 28040 31408
rect 27988 31365 27997 31399
rect 27997 31365 28031 31399
rect 28031 31365 28040 31399
rect 27988 31356 28040 31365
rect 17592 31331 17644 31340
rect 17592 31297 17601 31331
rect 17601 31297 17635 31331
rect 17635 31297 17644 31331
rect 17592 31288 17644 31297
rect 17684 31331 17736 31340
rect 17684 31297 17693 31331
rect 17693 31297 17727 31331
rect 17727 31297 17736 31331
rect 17684 31288 17736 31297
rect 17776 31331 17828 31340
rect 17776 31297 17785 31331
rect 17785 31297 17819 31331
rect 17819 31297 17828 31331
rect 17776 31288 17828 31297
rect 18052 31288 18104 31340
rect 18696 31288 18748 31340
rect 18788 31331 18840 31340
rect 18788 31297 18797 31331
rect 18797 31297 18831 31331
rect 18831 31297 18840 31331
rect 18788 31288 18840 31297
rect 19156 31288 19208 31340
rect 19708 31331 19760 31340
rect 19708 31297 19717 31331
rect 19717 31297 19751 31331
rect 19751 31297 19760 31331
rect 19708 31288 19760 31297
rect 20536 31331 20588 31340
rect 20536 31297 20545 31331
rect 20545 31297 20579 31331
rect 20579 31297 20588 31331
rect 20536 31288 20588 31297
rect 20628 31331 20680 31340
rect 20628 31297 20637 31331
rect 20637 31297 20671 31331
rect 20671 31297 20680 31331
rect 20628 31288 20680 31297
rect 20720 31288 20772 31340
rect 21088 31288 21140 31340
rect 21180 31263 21232 31272
rect 21180 31229 21189 31263
rect 21189 31229 21223 31263
rect 21223 31229 21232 31263
rect 21180 31220 21232 31229
rect 21640 31288 21692 31340
rect 21824 31331 21876 31340
rect 21824 31297 21833 31331
rect 21833 31297 21867 31331
rect 21867 31297 21876 31331
rect 21824 31288 21876 31297
rect 19524 31152 19576 31204
rect 21732 31220 21784 31272
rect 21456 31152 21508 31204
rect 21548 31152 21600 31204
rect 22560 31288 22612 31340
rect 22836 31331 22888 31340
rect 22836 31297 22845 31331
rect 22845 31297 22879 31331
rect 22879 31297 22888 31331
rect 22836 31288 22888 31297
rect 23020 31331 23072 31340
rect 23020 31297 23029 31331
rect 23029 31297 23063 31331
rect 23063 31297 23072 31331
rect 23020 31288 23072 31297
rect 23296 31331 23348 31340
rect 23296 31297 23305 31331
rect 23305 31297 23339 31331
rect 23339 31297 23348 31331
rect 23296 31288 23348 31297
rect 25412 31331 25464 31340
rect 25412 31297 25421 31331
rect 25421 31297 25455 31331
rect 25455 31297 25464 31331
rect 25412 31288 25464 31297
rect 25596 31331 25648 31340
rect 25596 31297 25605 31331
rect 25605 31297 25639 31331
rect 25639 31297 25648 31331
rect 25596 31288 25648 31297
rect 24584 31220 24636 31272
rect 26424 31288 26476 31340
rect 27160 31331 27212 31340
rect 27160 31297 27169 31331
rect 27169 31297 27203 31331
rect 27203 31297 27212 31331
rect 27160 31288 27212 31297
rect 26516 31220 26568 31272
rect 26792 31220 26844 31272
rect 17868 31084 17920 31136
rect 18328 31127 18380 31136
rect 18328 31093 18337 31127
rect 18337 31093 18371 31127
rect 18371 31093 18380 31127
rect 18328 31084 18380 31093
rect 19340 31084 19392 31136
rect 26700 31195 26752 31204
rect 26700 31161 26709 31195
rect 26709 31161 26743 31195
rect 26743 31161 26752 31195
rect 26700 31152 26752 31161
rect 27712 31263 27764 31272
rect 27712 31229 27721 31263
rect 27721 31229 27755 31263
rect 27755 31229 27764 31263
rect 27712 31220 27764 31229
rect 29644 31331 29696 31340
rect 29644 31297 29653 31331
rect 29653 31297 29687 31331
rect 29687 31297 29696 31331
rect 29644 31288 29696 31297
rect 29184 31152 29236 31204
rect 23020 31084 23072 31136
rect 25412 31084 25464 31136
rect 26424 31084 26476 31136
rect 27436 31084 27488 31136
rect 27712 31084 27764 31136
rect 29000 31084 29052 31136
rect 29552 31084 29604 31136
rect 31668 31288 31720 31340
rect 31944 31263 31996 31272
rect 31944 31229 31953 31263
rect 31953 31229 31987 31263
rect 31987 31229 31996 31263
rect 31944 31220 31996 31229
rect 34520 31331 34572 31340
rect 34520 31297 34529 31331
rect 34529 31297 34563 31331
rect 34563 31297 34572 31331
rect 34520 31288 34572 31297
rect 34152 31263 34204 31272
rect 34152 31229 34161 31263
rect 34161 31229 34195 31263
rect 34195 31229 34204 31263
rect 34152 31220 34204 31229
rect 35256 31220 35308 31272
rect 36544 31263 36596 31272
rect 36544 31229 36553 31263
rect 36553 31229 36587 31263
rect 36587 31229 36596 31263
rect 36544 31220 36596 31229
rect 32956 31084 33008 31136
rect 35992 31084 36044 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 6368 30880 6420 30932
rect 3976 30676 4028 30728
rect 5632 30719 5684 30728
rect 5632 30685 5641 30719
rect 5641 30685 5675 30719
rect 5675 30685 5684 30719
rect 5632 30676 5684 30685
rect 8392 30880 8444 30932
rect 8484 30880 8536 30932
rect 7472 30744 7524 30796
rect 9588 30880 9640 30932
rect 14464 30923 14516 30932
rect 14464 30889 14473 30923
rect 14473 30889 14507 30923
rect 14507 30889 14516 30923
rect 14464 30880 14516 30889
rect 16212 30880 16264 30932
rect 17592 30880 17644 30932
rect 11612 30812 11664 30864
rect 20996 30880 21048 30932
rect 21916 30880 21968 30932
rect 24400 30880 24452 30932
rect 25136 30880 25188 30932
rect 16856 30812 16908 30864
rect 17132 30812 17184 30864
rect 18052 30812 18104 30864
rect 20352 30855 20404 30864
rect 20352 30821 20361 30855
rect 20361 30821 20395 30855
rect 20395 30821 20404 30855
rect 20352 30812 20404 30821
rect 20720 30855 20772 30864
rect 20720 30821 20729 30855
rect 20729 30821 20763 30855
rect 20763 30821 20772 30855
rect 20720 30812 20772 30821
rect 22560 30812 22612 30864
rect 23296 30812 23348 30864
rect 9496 30787 9548 30796
rect 9496 30753 9505 30787
rect 9505 30753 9539 30787
rect 9539 30753 9548 30787
rect 9496 30744 9548 30753
rect 16948 30744 17000 30796
rect 24584 30787 24636 30796
rect 24584 30753 24593 30787
rect 24593 30753 24627 30787
rect 24627 30753 24636 30787
rect 27160 30880 27212 30932
rect 28264 30880 28316 30932
rect 29644 30880 29696 30932
rect 33324 30880 33376 30932
rect 24584 30744 24636 30753
rect 11704 30676 11756 30728
rect 4252 30540 4304 30592
rect 6184 30651 6236 30660
rect 6184 30617 6193 30651
rect 6193 30617 6227 30651
rect 6227 30617 6236 30651
rect 6184 30608 6236 30617
rect 9588 30608 9640 30660
rect 13268 30608 13320 30660
rect 13360 30608 13412 30660
rect 7840 30583 7892 30592
rect 7840 30549 7849 30583
rect 7849 30549 7883 30583
rect 7883 30549 7892 30583
rect 7840 30540 7892 30549
rect 8024 30540 8076 30592
rect 10232 30540 10284 30592
rect 13728 30651 13780 30660
rect 13728 30617 13737 30651
rect 13737 30617 13771 30651
rect 13771 30617 13780 30651
rect 13728 30608 13780 30617
rect 14464 30676 14516 30728
rect 14648 30719 14700 30728
rect 14648 30685 14657 30719
rect 14657 30685 14691 30719
rect 14691 30685 14700 30719
rect 14648 30676 14700 30685
rect 14740 30676 14792 30728
rect 16580 30719 16632 30728
rect 16580 30685 16589 30719
rect 16589 30685 16623 30719
rect 16623 30685 16632 30719
rect 16580 30676 16632 30685
rect 16672 30719 16724 30728
rect 16672 30685 16682 30719
rect 16682 30685 16716 30719
rect 16716 30685 16724 30719
rect 16672 30676 16724 30685
rect 16856 30719 16908 30728
rect 16856 30685 16865 30719
rect 16865 30685 16899 30719
rect 16899 30685 16908 30719
rect 16856 30676 16908 30685
rect 17408 30676 17460 30728
rect 17592 30676 17644 30728
rect 19064 30719 19116 30728
rect 19064 30685 19073 30719
rect 19073 30685 19107 30719
rect 19107 30685 19116 30719
rect 19064 30676 19116 30685
rect 19524 30719 19576 30728
rect 19524 30685 19533 30719
rect 19533 30685 19567 30719
rect 19567 30685 19576 30719
rect 19524 30676 19576 30685
rect 20260 30719 20312 30728
rect 20260 30685 20269 30719
rect 20269 30685 20303 30719
rect 20303 30685 20312 30719
rect 20260 30676 20312 30685
rect 20444 30676 20496 30728
rect 14096 30583 14148 30592
rect 14096 30549 14105 30583
rect 14105 30549 14139 30583
rect 14139 30549 14148 30583
rect 14096 30540 14148 30549
rect 14372 30540 14424 30592
rect 15936 30540 15988 30592
rect 16304 30540 16356 30592
rect 16672 30540 16724 30592
rect 18512 30608 18564 30660
rect 20352 30608 20404 30660
rect 21272 30676 21324 30728
rect 21364 30719 21416 30728
rect 21364 30685 21373 30719
rect 21373 30685 21407 30719
rect 21407 30685 21416 30719
rect 21364 30676 21416 30685
rect 25412 30676 25464 30728
rect 25964 30676 26016 30728
rect 26148 30719 26200 30728
rect 26148 30685 26157 30719
rect 26157 30685 26191 30719
rect 26191 30685 26200 30719
rect 26148 30676 26200 30685
rect 24584 30608 24636 30660
rect 26792 30744 26844 30796
rect 27620 30744 27672 30796
rect 28632 30787 28684 30796
rect 28632 30753 28641 30787
rect 28641 30753 28675 30787
rect 28675 30753 28684 30787
rect 28632 30744 28684 30753
rect 30656 30787 30708 30796
rect 30656 30753 30665 30787
rect 30665 30753 30699 30787
rect 30699 30753 30708 30787
rect 30656 30744 30708 30753
rect 31024 30744 31076 30796
rect 31668 30744 31720 30796
rect 26424 30719 26476 30728
rect 26424 30685 26433 30719
rect 26433 30685 26467 30719
rect 26467 30685 26476 30719
rect 26424 30676 26476 30685
rect 26608 30676 26660 30728
rect 27436 30676 27488 30728
rect 31944 30676 31996 30728
rect 32496 30676 32548 30728
rect 32772 30744 32824 30796
rect 33140 30787 33192 30796
rect 33140 30753 33149 30787
rect 33149 30753 33183 30787
rect 33183 30753 33192 30787
rect 33140 30744 33192 30753
rect 34152 30880 34204 30932
rect 35440 30923 35492 30932
rect 35440 30889 35449 30923
rect 35449 30889 35483 30923
rect 35483 30889 35492 30923
rect 35440 30880 35492 30889
rect 33968 30744 34020 30796
rect 17224 30583 17276 30592
rect 17224 30549 17233 30583
rect 17233 30549 17267 30583
rect 17267 30549 17276 30583
rect 17224 30540 17276 30549
rect 17960 30540 18012 30592
rect 18144 30540 18196 30592
rect 18788 30540 18840 30592
rect 19524 30540 19576 30592
rect 20076 30540 20128 30592
rect 20904 30583 20956 30592
rect 20904 30549 20913 30583
rect 20913 30549 20947 30583
rect 20947 30549 20956 30583
rect 20904 30540 20956 30549
rect 23572 30540 23624 30592
rect 29000 30608 29052 30660
rect 30932 30651 30984 30660
rect 30932 30617 30941 30651
rect 30941 30617 30975 30651
rect 30975 30617 30984 30651
rect 30932 30608 30984 30617
rect 33692 30608 33744 30660
rect 36544 30608 36596 30660
rect 28448 30583 28500 30592
rect 28448 30549 28457 30583
rect 28457 30549 28491 30583
rect 28491 30549 28500 30583
rect 28448 30540 28500 30549
rect 30840 30540 30892 30592
rect 31300 30540 31352 30592
rect 33324 30583 33376 30592
rect 33324 30549 33333 30583
rect 33333 30549 33367 30583
rect 33367 30549 33376 30583
rect 33324 30540 33376 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 5264 30268 5316 30320
rect 6184 30336 6236 30388
rect 4252 30175 4304 30184
rect 4252 30141 4261 30175
rect 4261 30141 4295 30175
rect 4295 30141 4304 30175
rect 4252 30132 4304 30141
rect 7656 30336 7708 30388
rect 7748 30336 7800 30388
rect 8024 30336 8076 30388
rect 9588 30336 9640 30388
rect 13452 30336 13504 30388
rect 15016 30336 15068 30388
rect 18052 30336 18104 30388
rect 19800 30336 19852 30388
rect 7288 30200 7340 30252
rect 7748 30243 7800 30252
rect 7748 30209 7757 30243
rect 7757 30209 7791 30243
rect 7791 30209 7800 30243
rect 7748 30200 7800 30209
rect 7932 30200 7984 30252
rect 9956 30268 10008 30320
rect 19524 30268 19576 30320
rect 8576 30243 8628 30252
rect 8576 30209 8585 30243
rect 8585 30209 8619 30243
rect 8619 30209 8628 30243
rect 8576 30200 8628 30209
rect 9496 30200 9548 30252
rect 10048 30200 10100 30252
rect 11520 30200 11572 30252
rect 11704 30243 11756 30252
rect 11704 30209 11714 30243
rect 11714 30209 11748 30243
rect 11748 30209 11756 30243
rect 11704 30200 11756 30209
rect 11888 30243 11940 30252
rect 11888 30209 11897 30243
rect 11897 30209 11931 30243
rect 11931 30209 11940 30243
rect 11888 30200 11940 30209
rect 12164 30200 12216 30252
rect 12348 30200 12400 30252
rect 13728 30200 13780 30252
rect 15200 30200 15252 30252
rect 16120 30200 16172 30252
rect 16488 30200 16540 30252
rect 15292 30132 15344 30184
rect 16672 30132 16724 30184
rect 16764 30132 16816 30184
rect 16948 30132 17000 30184
rect 17224 30132 17276 30184
rect 5264 29996 5316 30048
rect 5724 29996 5776 30048
rect 6828 29996 6880 30048
rect 9496 30064 9548 30116
rect 10692 30064 10744 30116
rect 7932 29996 7984 30048
rect 9404 29996 9456 30048
rect 12256 30039 12308 30048
rect 12256 30005 12265 30039
rect 12265 30005 12299 30039
rect 12299 30005 12308 30039
rect 12256 29996 12308 30005
rect 14556 30064 14608 30116
rect 15844 30064 15896 30116
rect 18512 30243 18564 30252
rect 18512 30209 18521 30243
rect 18521 30209 18555 30243
rect 18555 30209 18564 30243
rect 18512 30200 18564 30209
rect 18604 30243 18656 30252
rect 18604 30209 18613 30243
rect 18613 30209 18647 30243
rect 18647 30209 18656 30243
rect 18604 30200 18656 30209
rect 18328 30132 18380 30184
rect 18696 30132 18748 30184
rect 18972 30200 19024 30252
rect 19064 30200 19116 30252
rect 19984 30268 20036 30320
rect 20352 30336 20404 30388
rect 21088 30336 21140 30388
rect 23848 30336 23900 30388
rect 20628 30311 20680 30320
rect 20628 30277 20637 30311
rect 20637 30277 20671 30311
rect 20671 30277 20680 30311
rect 20628 30268 20680 30277
rect 21180 30268 21232 30320
rect 22652 30268 22704 30320
rect 23204 30268 23256 30320
rect 23388 30311 23440 30320
rect 23388 30277 23397 30311
rect 23397 30277 23431 30311
rect 23431 30277 23440 30311
rect 23388 30268 23440 30277
rect 24676 30268 24728 30320
rect 22008 30200 22060 30252
rect 22928 30200 22980 30252
rect 23112 30200 23164 30252
rect 26608 30268 26660 30320
rect 25780 30200 25832 30252
rect 25964 30243 26016 30252
rect 25964 30209 25973 30243
rect 25973 30209 26007 30243
rect 26007 30209 26016 30243
rect 25964 30200 26016 30209
rect 26148 30200 26200 30252
rect 26240 30200 26292 30252
rect 26516 30200 26568 30252
rect 29092 30379 29144 30388
rect 29092 30345 29101 30379
rect 29101 30345 29135 30379
rect 29135 30345 29144 30379
rect 29092 30336 29144 30345
rect 27804 30268 27856 30320
rect 30656 30268 30708 30320
rect 31024 30268 31076 30320
rect 29828 30200 29880 30252
rect 31300 30200 31352 30252
rect 27344 30132 27396 30184
rect 30840 30132 30892 30184
rect 32956 30336 33008 30388
rect 32036 30200 32088 30252
rect 32312 30243 32364 30252
rect 32312 30209 32321 30243
rect 32321 30209 32355 30243
rect 32355 30209 32364 30243
rect 32312 30200 32364 30209
rect 33048 30268 33100 30320
rect 33232 30268 33284 30320
rect 35992 30268 36044 30320
rect 32496 30243 32548 30252
rect 32496 30209 32505 30243
rect 32505 30209 32539 30243
rect 32539 30209 32548 30243
rect 32496 30200 32548 30209
rect 17408 29996 17460 30048
rect 17868 30039 17920 30048
rect 17868 30005 17877 30039
rect 17877 30005 17911 30039
rect 17911 30005 17920 30039
rect 17868 29996 17920 30005
rect 18328 29996 18380 30048
rect 20352 30064 20404 30116
rect 18696 29996 18748 30048
rect 19892 29996 19944 30048
rect 20444 29996 20496 30048
rect 20536 29996 20588 30048
rect 21548 30064 21600 30116
rect 22284 30064 22336 30116
rect 26056 30064 26108 30116
rect 26608 30064 26660 30116
rect 27804 30064 27856 30116
rect 27988 30064 28040 30116
rect 33324 30064 33376 30116
rect 20812 30039 20864 30048
rect 20812 30005 20821 30039
rect 20821 30005 20855 30039
rect 20855 30005 20864 30039
rect 20812 29996 20864 30005
rect 23940 29996 23992 30048
rect 25320 29996 25372 30048
rect 25780 29996 25832 30048
rect 26700 29996 26752 30048
rect 29920 29996 29972 30048
rect 30564 29996 30616 30048
rect 32956 29996 33008 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 10692 29835 10744 29844
rect 10692 29801 10701 29835
rect 10701 29801 10735 29835
rect 10735 29801 10744 29835
rect 10692 29792 10744 29801
rect 12256 29792 12308 29844
rect 3976 29588 4028 29640
rect 6920 29724 6972 29776
rect 6828 29656 6880 29708
rect 12624 29792 12676 29844
rect 16580 29792 16632 29844
rect 17408 29792 17460 29844
rect 15292 29724 15344 29776
rect 18328 29724 18380 29776
rect 18696 29724 18748 29776
rect 18880 29767 18932 29776
rect 18880 29733 18889 29767
rect 18889 29733 18923 29767
rect 18923 29733 18932 29767
rect 18880 29724 18932 29733
rect 19800 29792 19852 29844
rect 20076 29792 20128 29844
rect 20720 29792 20772 29844
rect 21272 29792 21324 29844
rect 22008 29792 22060 29844
rect 24124 29792 24176 29844
rect 24400 29792 24452 29844
rect 20628 29767 20680 29776
rect 20628 29733 20637 29767
rect 20637 29733 20671 29767
rect 20671 29733 20680 29767
rect 20628 29724 20680 29733
rect 8300 29631 8352 29640
rect 8300 29597 8309 29631
rect 8309 29597 8343 29631
rect 8343 29597 8352 29631
rect 8300 29588 8352 29597
rect 4068 29495 4120 29504
rect 4068 29461 4077 29495
rect 4077 29461 4111 29495
rect 4111 29461 4120 29495
rect 4068 29452 4120 29461
rect 5448 29495 5500 29504
rect 5448 29461 5457 29495
rect 5457 29461 5491 29495
rect 5491 29461 5500 29495
rect 5448 29452 5500 29461
rect 6092 29520 6144 29572
rect 8392 29520 8444 29572
rect 6828 29452 6880 29504
rect 12716 29631 12768 29640
rect 12716 29597 12725 29631
rect 12725 29597 12759 29631
rect 12759 29597 12768 29631
rect 12716 29588 12768 29597
rect 9680 29520 9732 29572
rect 13544 29631 13596 29640
rect 13544 29597 13553 29631
rect 13553 29597 13587 29631
rect 13587 29597 13596 29631
rect 13544 29588 13596 29597
rect 13912 29588 13964 29640
rect 14096 29588 14148 29640
rect 15108 29588 15160 29640
rect 15476 29631 15528 29640
rect 15476 29597 15485 29631
rect 15485 29597 15519 29631
rect 15519 29597 15528 29631
rect 15476 29588 15528 29597
rect 15660 29631 15712 29640
rect 15660 29597 15669 29631
rect 15669 29597 15703 29631
rect 15703 29597 15712 29631
rect 15660 29588 15712 29597
rect 15844 29588 15896 29640
rect 18052 29656 18104 29708
rect 16120 29631 16172 29640
rect 16120 29597 16129 29631
rect 16129 29597 16163 29631
rect 16163 29597 16172 29631
rect 16120 29588 16172 29597
rect 9036 29452 9088 29504
rect 9956 29452 10008 29504
rect 13268 29495 13320 29504
rect 13268 29461 13277 29495
rect 13277 29461 13311 29495
rect 13311 29461 13320 29495
rect 13268 29452 13320 29461
rect 15016 29520 15068 29572
rect 16028 29563 16080 29572
rect 16028 29529 16037 29563
rect 16037 29529 16071 29563
rect 16071 29529 16080 29563
rect 16028 29520 16080 29529
rect 16396 29520 16448 29572
rect 18144 29588 18196 29640
rect 18512 29631 18564 29640
rect 18512 29597 18521 29631
rect 18521 29597 18555 29631
rect 18555 29597 18564 29631
rect 18512 29588 18564 29597
rect 18972 29656 19024 29708
rect 19708 29656 19760 29708
rect 19892 29656 19944 29708
rect 18696 29631 18748 29640
rect 18696 29597 18705 29631
rect 18705 29597 18739 29631
rect 18739 29597 18748 29631
rect 18696 29588 18748 29597
rect 19156 29588 19208 29640
rect 20536 29588 20588 29640
rect 21640 29656 21692 29708
rect 21272 29588 21324 29640
rect 21456 29588 21508 29640
rect 16764 29452 16816 29504
rect 16856 29495 16908 29504
rect 16856 29461 16865 29495
rect 16865 29461 16899 29495
rect 16899 29461 16908 29495
rect 16856 29452 16908 29461
rect 16948 29495 17000 29504
rect 16948 29461 16957 29495
rect 16957 29461 16991 29495
rect 16991 29461 17000 29495
rect 16948 29452 17000 29461
rect 17040 29495 17092 29504
rect 17040 29461 17049 29495
rect 17049 29461 17083 29495
rect 17083 29461 17092 29495
rect 17040 29452 17092 29461
rect 22284 29520 22336 29572
rect 22744 29588 22796 29640
rect 22928 29631 22980 29640
rect 22928 29597 22932 29631
rect 22932 29597 22966 29631
rect 22966 29597 22980 29631
rect 22928 29588 22980 29597
rect 23848 29724 23900 29776
rect 23480 29656 23532 29708
rect 23204 29631 23256 29640
rect 23204 29597 23249 29631
rect 23249 29597 23256 29631
rect 23204 29588 23256 29597
rect 23388 29631 23440 29640
rect 23388 29597 23397 29631
rect 23397 29597 23431 29631
rect 23431 29597 23440 29631
rect 23388 29588 23440 29597
rect 23756 29631 23808 29640
rect 23756 29597 23765 29631
rect 23765 29597 23799 29631
rect 23799 29597 23808 29631
rect 23756 29588 23808 29597
rect 25136 29724 25188 29776
rect 24584 29656 24636 29708
rect 24676 29699 24728 29708
rect 24676 29665 24685 29699
rect 24685 29665 24719 29699
rect 24719 29665 24728 29699
rect 24676 29656 24728 29665
rect 24308 29588 24360 29640
rect 24952 29588 25004 29640
rect 26056 29724 26108 29776
rect 26056 29588 26108 29640
rect 26332 29588 26384 29640
rect 26424 29631 26476 29640
rect 26424 29597 26433 29631
rect 26433 29597 26467 29631
rect 26467 29597 26476 29631
rect 26424 29588 26476 29597
rect 26700 29724 26752 29776
rect 27344 29724 27396 29776
rect 28724 29724 28776 29776
rect 29276 29724 29328 29776
rect 30380 29724 30432 29776
rect 26792 29631 26844 29640
rect 26792 29597 26801 29631
rect 26801 29597 26835 29631
rect 26835 29597 26844 29631
rect 26792 29588 26844 29597
rect 27344 29631 27396 29640
rect 27344 29597 27353 29631
rect 27353 29597 27387 29631
rect 27387 29597 27396 29631
rect 27344 29588 27396 29597
rect 27620 29699 27672 29708
rect 27620 29665 27629 29699
rect 27629 29665 27663 29699
rect 27663 29665 27672 29699
rect 27620 29656 27672 29665
rect 20996 29452 21048 29504
rect 21824 29452 21876 29504
rect 22652 29452 22704 29504
rect 23296 29452 23348 29504
rect 23572 29495 23624 29504
rect 23572 29461 23581 29495
rect 23581 29461 23615 29495
rect 23615 29461 23624 29495
rect 23572 29452 23624 29461
rect 25780 29452 25832 29504
rect 26516 29452 26568 29504
rect 29000 29656 29052 29708
rect 27988 29452 28040 29504
rect 28724 29588 28776 29640
rect 29644 29588 29696 29640
rect 29828 29631 29880 29640
rect 29828 29597 29837 29631
rect 29837 29597 29871 29631
rect 29871 29597 29880 29631
rect 29828 29588 29880 29597
rect 28356 29495 28408 29504
rect 28356 29461 28365 29495
rect 28365 29461 28399 29495
rect 28399 29461 28408 29495
rect 28356 29452 28408 29461
rect 29276 29495 29328 29504
rect 29276 29461 29285 29495
rect 29285 29461 29319 29495
rect 29319 29461 29328 29495
rect 29276 29452 29328 29461
rect 29552 29495 29604 29504
rect 29552 29461 29561 29495
rect 29561 29461 29595 29495
rect 29595 29461 29604 29495
rect 29552 29452 29604 29461
rect 29828 29452 29880 29504
rect 30012 29631 30064 29640
rect 30012 29597 30021 29631
rect 30021 29597 30055 29631
rect 30055 29597 30064 29631
rect 30012 29588 30064 29597
rect 30196 29631 30248 29640
rect 30196 29597 30205 29631
rect 30205 29597 30239 29631
rect 30239 29597 30248 29631
rect 30196 29588 30248 29597
rect 34060 29724 34112 29776
rect 34244 29724 34296 29776
rect 30564 29631 30616 29640
rect 30564 29597 30573 29631
rect 30573 29597 30607 29631
rect 30607 29597 30616 29631
rect 30564 29588 30616 29597
rect 30748 29588 30800 29640
rect 31024 29588 31076 29640
rect 31300 29588 31352 29640
rect 31668 29588 31720 29640
rect 34796 29631 34848 29640
rect 34796 29597 34805 29631
rect 34805 29597 34839 29631
rect 34839 29597 34848 29631
rect 34796 29588 34848 29597
rect 30656 29563 30708 29572
rect 30656 29529 30665 29563
rect 30665 29529 30699 29563
rect 30699 29529 30708 29563
rect 30656 29520 30708 29529
rect 31116 29520 31168 29572
rect 34336 29520 34388 29572
rect 34980 29520 35032 29572
rect 30932 29495 30984 29504
rect 30932 29461 30941 29495
rect 30941 29461 30975 29495
rect 30975 29461 30984 29495
rect 30932 29452 30984 29461
rect 33324 29452 33376 29504
rect 34520 29495 34572 29504
rect 34520 29461 34529 29495
rect 34529 29461 34563 29495
rect 34563 29461 34572 29495
rect 34520 29452 34572 29461
rect 35992 29452 36044 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4068 29248 4120 29300
rect 6828 29248 6880 29300
rect 6092 29180 6144 29232
rect 8300 29248 8352 29300
rect 10692 29248 10744 29300
rect 16764 29248 16816 29300
rect 5264 29112 5316 29164
rect 7012 29044 7064 29096
rect 7932 29112 7984 29164
rect 6920 28976 6972 29028
rect 17960 29180 18012 29232
rect 18696 29248 18748 29300
rect 18972 29248 19024 29300
rect 12716 29112 12768 29164
rect 16672 29112 16724 29164
rect 16856 29112 16908 29164
rect 17224 29112 17276 29164
rect 17500 29112 17552 29164
rect 17684 29112 17736 29164
rect 18420 29112 18472 29164
rect 18604 29112 18656 29164
rect 9128 29044 9180 29096
rect 10968 29044 11020 29096
rect 16028 29044 16080 29096
rect 20352 29180 20404 29232
rect 20904 29223 20956 29232
rect 20904 29189 20913 29223
rect 20913 29189 20947 29223
rect 20947 29189 20956 29223
rect 20904 29180 20956 29189
rect 19892 29112 19944 29164
rect 20628 29112 20680 29164
rect 21456 29248 21508 29300
rect 21640 29248 21692 29300
rect 21088 29155 21140 29164
rect 21088 29121 21097 29155
rect 21097 29121 21131 29155
rect 21131 29121 21140 29155
rect 21088 29112 21140 29121
rect 21640 29112 21692 29164
rect 21824 29155 21876 29164
rect 21824 29121 21833 29155
rect 21833 29121 21867 29155
rect 21867 29121 21876 29155
rect 21824 29112 21876 29121
rect 22008 29155 22060 29164
rect 22008 29121 22015 29155
rect 22015 29121 22060 29155
rect 22008 29112 22060 29121
rect 22100 29155 22152 29164
rect 22100 29121 22109 29155
rect 22109 29121 22143 29155
rect 22143 29121 22152 29155
rect 22100 29112 22152 29121
rect 22192 29155 22244 29164
rect 22192 29121 22201 29155
rect 22201 29121 22235 29155
rect 22235 29121 22244 29155
rect 22192 29112 22244 29121
rect 22376 29180 22428 29232
rect 23204 29180 23256 29232
rect 22560 29155 22612 29164
rect 22560 29121 22569 29155
rect 22569 29121 22603 29155
rect 22603 29121 22612 29155
rect 22560 29112 22612 29121
rect 22652 29112 22704 29164
rect 23020 29155 23072 29164
rect 23020 29121 23029 29155
rect 23029 29121 23063 29155
rect 23063 29121 23072 29155
rect 23020 29112 23072 29121
rect 23664 29223 23716 29232
rect 23664 29189 23673 29223
rect 23673 29189 23707 29223
rect 23707 29189 23716 29223
rect 23664 29180 23716 29189
rect 23848 29248 23900 29300
rect 23940 29112 23992 29164
rect 25412 29112 25464 29164
rect 12900 29019 12952 29028
rect 12900 28985 12909 29019
rect 12909 28985 12943 29019
rect 12943 28985 12952 29019
rect 12900 28976 12952 28985
rect 13728 28976 13780 29028
rect 4620 28908 4672 28960
rect 5356 28908 5408 28960
rect 6552 28908 6604 28960
rect 8392 28908 8444 28960
rect 8484 28908 8536 28960
rect 18420 28908 18472 28960
rect 18604 28951 18656 28960
rect 18604 28917 18613 28951
rect 18613 28917 18647 28951
rect 18647 28917 18656 28951
rect 18604 28908 18656 28917
rect 19156 28908 19208 28960
rect 19892 28908 19944 28960
rect 21272 28954 21324 29006
rect 23204 28951 23256 28960
rect 23204 28917 23213 28951
rect 23213 28917 23247 28951
rect 23247 28917 23256 28951
rect 23204 28908 23256 28917
rect 23940 28976 23992 29028
rect 25596 29155 25648 29164
rect 25596 29121 25605 29155
rect 25605 29121 25639 29155
rect 25639 29121 25648 29155
rect 25596 29112 25648 29121
rect 26424 29248 26476 29300
rect 26516 29248 26568 29300
rect 27344 29248 27396 29300
rect 25964 29112 26016 29164
rect 26884 29112 26936 29164
rect 28356 29248 28408 29300
rect 29000 29291 29052 29300
rect 29000 29257 29009 29291
rect 29009 29257 29043 29291
rect 29043 29257 29052 29291
rect 29000 29248 29052 29257
rect 29276 29248 29328 29300
rect 30932 29248 30984 29300
rect 31576 29291 31628 29300
rect 31576 29257 31585 29291
rect 31585 29257 31619 29291
rect 31619 29257 31628 29291
rect 31576 29248 31628 29257
rect 31668 29248 31720 29300
rect 28632 29112 28684 29164
rect 30840 29180 30892 29232
rect 31484 29155 31536 29164
rect 31484 29121 31493 29155
rect 31493 29121 31527 29155
rect 31527 29121 31536 29155
rect 31484 29112 31536 29121
rect 34796 29248 34848 29300
rect 34336 29180 34388 29232
rect 32312 29155 32364 29164
rect 32312 29121 32321 29155
rect 32321 29121 32355 29155
rect 32355 29121 32364 29155
rect 32312 29112 32364 29121
rect 30012 29044 30064 29096
rect 33048 29155 33100 29164
rect 33048 29121 33057 29155
rect 33057 29121 33091 29155
rect 33091 29121 33100 29155
rect 33048 29112 33100 29121
rect 34520 29112 34572 29164
rect 34980 29112 35032 29164
rect 36636 29155 36688 29164
rect 36636 29121 36645 29155
rect 36645 29121 36679 29155
rect 36679 29121 36688 29155
rect 36636 29112 36688 29121
rect 36820 29155 36872 29164
rect 36820 29121 36829 29155
rect 36829 29121 36863 29155
rect 36863 29121 36872 29155
rect 36820 29112 36872 29121
rect 26700 28976 26752 29028
rect 27068 28976 27120 29028
rect 24032 28951 24084 28960
rect 24032 28917 24041 28951
rect 24041 28917 24075 28951
rect 24075 28917 24084 28951
rect 24032 28908 24084 28917
rect 25412 28908 25464 28960
rect 25964 28908 26016 28960
rect 29276 28908 29328 28960
rect 30196 28908 30248 28960
rect 31116 28976 31168 29028
rect 33232 29044 33284 29096
rect 34704 28976 34756 29028
rect 37280 28976 37332 29028
rect 32404 28908 32456 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4620 28704 4672 28756
rect 8484 28704 8536 28756
rect 6552 28568 6604 28620
rect 20260 28704 20312 28756
rect 25596 28704 25648 28756
rect 16304 28636 16356 28688
rect 29092 28704 29144 28756
rect 29276 28747 29328 28756
rect 29276 28713 29285 28747
rect 29285 28713 29319 28747
rect 29319 28713 29328 28747
rect 29276 28704 29328 28713
rect 5448 28500 5500 28552
rect 5632 28500 5684 28552
rect 18328 28568 18380 28620
rect 18972 28568 19024 28620
rect 19616 28568 19668 28620
rect 4252 28407 4304 28416
rect 4252 28373 4261 28407
rect 4261 28373 4295 28407
rect 4295 28373 4304 28407
rect 4252 28364 4304 28373
rect 7196 28432 7248 28484
rect 8116 28432 8168 28484
rect 9956 28543 10008 28552
rect 9956 28509 9965 28543
rect 9965 28509 9999 28543
rect 9999 28509 10008 28543
rect 9956 28500 10008 28509
rect 13452 28500 13504 28552
rect 14280 28500 14332 28552
rect 16120 28543 16172 28552
rect 16120 28509 16129 28543
rect 16129 28509 16163 28543
rect 16163 28509 16172 28543
rect 16120 28500 16172 28509
rect 16212 28500 16264 28552
rect 16488 28543 16540 28552
rect 16488 28509 16497 28543
rect 16497 28509 16531 28543
rect 16531 28509 16540 28543
rect 16488 28500 16540 28509
rect 17960 28500 18012 28552
rect 19892 28568 19944 28620
rect 24492 28568 24544 28620
rect 10416 28432 10468 28484
rect 10508 28475 10560 28484
rect 10508 28441 10517 28475
rect 10517 28441 10551 28475
rect 10551 28441 10560 28475
rect 10508 28432 10560 28441
rect 11060 28432 11112 28484
rect 14096 28432 14148 28484
rect 16856 28432 16908 28484
rect 17868 28432 17920 28484
rect 19340 28432 19392 28484
rect 20628 28500 20680 28552
rect 20812 28543 20864 28552
rect 20812 28509 20821 28543
rect 20821 28509 20855 28543
rect 20855 28509 20864 28543
rect 20812 28500 20864 28509
rect 20996 28500 21048 28552
rect 21272 28500 21324 28552
rect 21640 28500 21692 28552
rect 22008 28500 22060 28552
rect 22376 28500 22428 28552
rect 22560 28500 22612 28552
rect 22928 28500 22980 28552
rect 23756 28500 23808 28552
rect 24676 28543 24728 28552
rect 24676 28509 24685 28543
rect 24685 28509 24719 28543
rect 24719 28509 24728 28543
rect 24676 28500 24728 28509
rect 24952 28543 25004 28552
rect 24952 28509 24961 28543
rect 24961 28509 24995 28543
rect 24995 28509 25004 28543
rect 24952 28500 25004 28509
rect 25320 28500 25372 28552
rect 25596 28500 25648 28552
rect 26148 28568 26200 28620
rect 30012 28611 30064 28620
rect 30012 28577 30021 28611
rect 30021 28577 30055 28611
rect 30055 28577 30064 28611
rect 30012 28568 30064 28577
rect 30104 28611 30156 28620
rect 30104 28577 30113 28611
rect 30113 28577 30147 28611
rect 30147 28577 30156 28611
rect 30104 28568 30156 28577
rect 31576 28636 31628 28688
rect 7932 28364 7984 28416
rect 11980 28407 12032 28416
rect 11980 28373 11989 28407
rect 11989 28373 12023 28407
rect 12023 28373 12032 28407
rect 11980 28364 12032 28373
rect 16488 28364 16540 28416
rect 19432 28364 19484 28416
rect 20168 28364 20220 28416
rect 21088 28364 21140 28416
rect 21548 28364 21600 28416
rect 23756 28364 23808 28416
rect 24400 28407 24452 28416
rect 24400 28373 24409 28407
rect 24409 28373 24443 28407
rect 24443 28373 24452 28407
rect 24400 28364 24452 28373
rect 24768 28475 24820 28484
rect 24768 28441 24777 28475
rect 24777 28441 24811 28475
rect 24811 28441 24820 28475
rect 24768 28432 24820 28441
rect 25872 28432 25924 28484
rect 24952 28364 25004 28416
rect 30380 28543 30432 28552
rect 30380 28509 30389 28543
rect 30389 28509 30423 28543
rect 30423 28509 30432 28543
rect 30380 28500 30432 28509
rect 30656 28475 30708 28484
rect 30656 28441 30665 28475
rect 30665 28441 30699 28475
rect 30699 28441 30708 28475
rect 30656 28432 30708 28441
rect 30196 28364 30248 28416
rect 30932 28364 30984 28416
rect 31484 28500 31536 28552
rect 32404 28568 32456 28620
rect 33324 28568 33376 28620
rect 33968 28568 34020 28620
rect 31760 28543 31812 28552
rect 31760 28509 31769 28543
rect 31769 28509 31803 28543
rect 31803 28509 31812 28543
rect 31760 28500 31812 28509
rect 34704 28543 34756 28552
rect 34704 28509 34713 28543
rect 34713 28509 34747 28543
rect 34747 28509 34756 28543
rect 34704 28500 34756 28509
rect 31944 28432 31996 28484
rect 34060 28432 34112 28484
rect 34428 28432 34480 28484
rect 35992 28432 36044 28484
rect 31116 28407 31168 28416
rect 31116 28373 31125 28407
rect 31125 28373 31159 28407
rect 31159 28373 31168 28407
rect 31116 28364 31168 28373
rect 31484 28407 31536 28416
rect 31484 28373 31493 28407
rect 31493 28373 31527 28407
rect 31527 28373 31536 28407
rect 31484 28364 31536 28373
rect 34152 28407 34204 28416
rect 34152 28373 34161 28407
rect 34161 28373 34195 28407
rect 34195 28373 34204 28407
rect 34152 28364 34204 28373
rect 34520 28407 34572 28416
rect 34520 28373 34529 28407
rect 34529 28373 34563 28407
rect 34563 28373 34572 28407
rect 34520 28364 34572 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4252 28160 4304 28212
rect 6828 28203 6880 28212
rect 6828 28169 6837 28203
rect 6837 28169 6871 28203
rect 6871 28169 6880 28203
rect 6828 28160 6880 28169
rect 4620 28092 4672 28144
rect 7196 28092 7248 28144
rect 5356 28024 5408 28076
rect 6000 28024 6052 28076
rect 7932 28092 7984 28144
rect 9680 28160 9732 28212
rect 10508 28160 10560 28212
rect 7472 27956 7524 28008
rect 6368 27863 6420 27872
rect 6368 27829 6377 27863
rect 6377 27829 6411 27863
rect 6411 27829 6420 27863
rect 6368 27820 6420 27829
rect 9772 28024 9824 28076
rect 8300 27956 8352 28008
rect 10140 27999 10192 28008
rect 10140 27965 10149 27999
rect 10149 27965 10183 27999
rect 10183 27965 10192 27999
rect 10140 27956 10192 27965
rect 11980 28160 12032 28212
rect 12532 28160 12584 28212
rect 13452 28160 13504 28212
rect 14004 28160 14056 28212
rect 16120 28160 16172 28212
rect 16580 28160 16632 28212
rect 15844 28092 15896 28144
rect 16856 28092 16908 28144
rect 11980 27999 12032 28008
rect 11980 27965 11989 27999
rect 11989 27965 12023 27999
rect 12023 27965 12032 27999
rect 11980 27956 12032 27965
rect 12072 27999 12124 28008
rect 12072 27965 12081 27999
rect 12081 27965 12115 27999
rect 12115 27965 12124 27999
rect 12072 27956 12124 27965
rect 13176 28024 13228 28076
rect 14372 28024 14424 28076
rect 14556 28024 14608 28076
rect 15200 28024 15252 28076
rect 16028 28024 16080 28076
rect 16764 28067 16816 28076
rect 16764 28033 16774 28067
rect 16774 28033 16808 28067
rect 16808 28033 16816 28067
rect 16764 28024 16816 28033
rect 17316 28024 17368 28076
rect 17868 28024 17920 28076
rect 18420 28160 18472 28212
rect 18788 28160 18840 28212
rect 18788 28024 18840 28076
rect 19156 28092 19208 28144
rect 20720 28092 20772 28144
rect 19340 27956 19392 28008
rect 19524 27956 19576 28008
rect 19892 28033 19911 28042
rect 19911 28033 19944 28042
rect 19892 27990 19944 28033
rect 20076 28067 20128 28076
rect 20076 28033 20085 28067
rect 20085 28033 20119 28067
rect 20119 28033 20128 28067
rect 20076 28024 20128 28033
rect 14648 27931 14700 27940
rect 14648 27897 14657 27931
rect 14657 27897 14691 27931
rect 14691 27897 14700 27931
rect 14648 27888 14700 27897
rect 15752 27888 15804 27940
rect 9496 27820 9548 27872
rect 9680 27820 9732 27872
rect 10968 27820 11020 27872
rect 12072 27820 12124 27872
rect 13636 27820 13688 27872
rect 14188 27863 14240 27872
rect 14188 27829 14197 27863
rect 14197 27829 14231 27863
rect 14231 27829 14240 27863
rect 14188 27820 14240 27829
rect 14464 27863 14516 27872
rect 14464 27829 14473 27863
rect 14473 27829 14507 27863
rect 14507 27829 14516 27863
rect 14464 27820 14516 27829
rect 15476 27820 15528 27872
rect 16120 27820 16172 27872
rect 17316 27863 17368 27872
rect 17316 27829 17325 27863
rect 17325 27829 17359 27863
rect 17359 27829 17368 27863
rect 17316 27820 17368 27829
rect 17408 27820 17460 27872
rect 17684 27820 17736 27872
rect 18236 27820 18288 27872
rect 19616 27888 19668 27940
rect 20352 27999 20404 28008
rect 20352 27965 20361 27999
rect 20361 27965 20395 27999
rect 20395 27965 20404 27999
rect 20352 27956 20404 27965
rect 19892 27820 19944 27872
rect 20536 27820 20588 27872
rect 23020 28160 23072 28212
rect 23296 28160 23348 28212
rect 24216 28160 24268 28212
rect 26792 28160 26844 28212
rect 29092 28160 29144 28212
rect 31484 28160 31536 28212
rect 31760 28160 31812 28212
rect 31944 28160 31996 28212
rect 33048 28160 33100 28212
rect 34428 28203 34480 28212
rect 34428 28169 34437 28203
rect 34437 28169 34471 28203
rect 34471 28169 34480 28203
rect 34428 28160 34480 28169
rect 34612 28160 34664 28212
rect 34704 28160 34756 28212
rect 37280 28160 37332 28212
rect 22192 28092 22244 28144
rect 21456 28024 21508 28076
rect 21640 28024 21692 28076
rect 23204 28024 23256 28076
rect 21824 27956 21876 28008
rect 21916 27999 21968 28008
rect 21916 27965 21925 27999
rect 21925 27965 21959 27999
rect 21959 27965 21968 27999
rect 21916 27956 21968 27965
rect 22928 27956 22980 28008
rect 23388 28067 23440 28076
rect 23388 28033 23397 28067
rect 23397 28033 23431 28067
rect 23431 28033 23440 28067
rect 23388 28024 23440 28033
rect 23572 28024 23624 28076
rect 23756 28067 23808 28076
rect 23756 28033 23765 28067
rect 23765 28033 23799 28067
rect 23799 28033 23808 28067
rect 23756 28024 23808 28033
rect 24032 28024 24084 28076
rect 24400 28024 24452 28076
rect 24676 28024 24728 28076
rect 21272 27820 21324 27872
rect 22284 27820 22336 27872
rect 30196 27956 30248 28008
rect 34152 28024 34204 28076
rect 34520 28024 34572 28076
rect 33140 27956 33192 28008
rect 33876 27956 33928 28008
rect 24216 27863 24268 27872
rect 24216 27829 24225 27863
rect 24225 27829 24259 27863
rect 24259 27829 24268 27863
rect 24216 27820 24268 27829
rect 24492 27863 24544 27872
rect 24492 27829 24501 27863
rect 24501 27829 24535 27863
rect 24535 27829 24544 27863
rect 24492 27820 24544 27829
rect 26516 27820 26568 27872
rect 28264 27820 28316 27872
rect 28816 27820 28868 27872
rect 29736 27820 29788 27872
rect 37556 27863 37608 27872
rect 37556 27829 37565 27863
rect 37565 27829 37599 27863
rect 37599 27829 37608 27863
rect 37556 27820 37608 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4620 27659 4672 27668
rect 4620 27625 4629 27659
rect 4629 27625 4663 27659
rect 4663 27625 4672 27659
rect 4620 27616 4672 27625
rect 8300 27659 8352 27668
rect 8300 27625 8309 27659
rect 8309 27625 8343 27659
rect 8343 27625 8352 27659
rect 8300 27616 8352 27625
rect 9496 27616 9548 27668
rect 9680 27616 9732 27668
rect 6368 27412 6420 27464
rect 6920 27455 6972 27464
rect 6920 27421 6929 27455
rect 6929 27421 6963 27455
rect 6963 27421 6972 27455
rect 9588 27548 9640 27600
rect 14096 27591 14148 27600
rect 14096 27557 14105 27591
rect 14105 27557 14139 27591
rect 14139 27557 14148 27591
rect 14096 27548 14148 27557
rect 14648 27659 14700 27668
rect 14648 27625 14657 27659
rect 14657 27625 14691 27659
rect 14691 27625 14700 27659
rect 14648 27616 14700 27625
rect 16028 27659 16080 27668
rect 16028 27625 16037 27659
rect 16037 27625 16071 27659
rect 16071 27625 16080 27659
rect 16028 27616 16080 27625
rect 20444 27616 20496 27668
rect 11980 27480 12032 27532
rect 6920 27412 6972 27421
rect 11060 27412 11112 27464
rect 10048 27387 10100 27396
rect 10048 27353 10057 27387
rect 10057 27353 10091 27387
rect 10091 27353 10100 27387
rect 10048 27344 10100 27353
rect 13728 27480 13780 27532
rect 13176 27412 13228 27464
rect 13544 27412 13596 27464
rect 13820 27412 13872 27464
rect 15568 27455 15620 27464
rect 15568 27421 15577 27455
rect 15577 27421 15611 27455
rect 15611 27421 15620 27455
rect 15568 27412 15620 27421
rect 6828 27319 6880 27328
rect 6828 27285 6837 27319
rect 6837 27285 6871 27319
rect 6871 27285 6880 27319
rect 6828 27276 6880 27285
rect 7564 27276 7616 27328
rect 11612 27319 11664 27328
rect 11612 27285 11621 27319
rect 11621 27285 11655 27319
rect 11655 27285 11664 27319
rect 11612 27276 11664 27285
rect 12532 27344 12584 27396
rect 14464 27387 14516 27396
rect 14464 27353 14473 27387
rect 14473 27353 14507 27387
rect 14507 27353 14516 27387
rect 14464 27344 14516 27353
rect 16120 27412 16172 27464
rect 16580 27412 16632 27464
rect 16672 27455 16724 27464
rect 16672 27421 16681 27455
rect 16681 27421 16715 27455
rect 16715 27421 16724 27455
rect 16672 27412 16724 27421
rect 16764 27455 16816 27464
rect 16764 27421 16774 27455
rect 16774 27421 16808 27455
rect 16808 27421 16816 27455
rect 16764 27412 16816 27421
rect 17132 27548 17184 27600
rect 17592 27548 17644 27600
rect 17684 27548 17736 27600
rect 18972 27548 19024 27600
rect 20168 27548 20220 27600
rect 20628 27548 20680 27600
rect 17868 27480 17920 27532
rect 18052 27480 18104 27532
rect 17408 27455 17460 27464
rect 17408 27421 17439 27455
rect 17439 27421 17460 27455
rect 17408 27412 17460 27421
rect 17500 27412 17552 27464
rect 17684 27455 17736 27464
rect 17684 27421 17693 27455
rect 17693 27421 17727 27455
rect 17727 27421 17736 27455
rect 17684 27412 17736 27421
rect 18144 27455 18196 27464
rect 18144 27421 18153 27455
rect 18153 27421 18187 27455
rect 18187 27421 18196 27455
rect 18144 27412 18196 27421
rect 21272 27480 21324 27532
rect 21732 27480 21784 27532
rect 18604 27455 18656 27464
rect 18604 27421 18613 27455
rect 18613 27421 18647 27455
rect 18647 27421 18656 27455
rect 18604 27412 18656 27421
rect 19340 27412 19392 27464
rect 23388 27616 23440 27668
rect 24216 27616 24268 27668
rect 12348 27276 12400 27328
rect 14280 27319 14332 27328
rect 14280 27285 14289 27319
rect 14289 27285 14323 27319
rect 14323 27285 14332 27319
rect 14280 27276 14332 27285
rect 14372 27319 14424 27328
rect 14372 27285 14381 27319
rect 14381 27285 14415 27319
rect 14415 27285 14424 27319
rect 14372 27276 14424 27285
rect 14556 27276 14608 27328
rect 15568 27276 15620 27328
rect 16856 27276 16908 27328
rect 18512 27387 18564 27396
rect 18512 27353 18521 27387
rect 18521 27353 18555 27387
rect 18555 27353 18564 27387
rect 18512 27344 18564 27353
rect 17776 27276 17828 27328
rect 18420 27276 18472 27328
rect 19432 27344 19484 27396
rect 19892 27344 19944 27396
rect 21088 27344 21140 27396
rect 21456 27344 21508 27396
rect 18788 27319 18840 27328
rect 18788 27285 18797 27319
rect 18797 27285 18831 27319
rect 18831 27285 18840 27319
rect 18788 27276 18840 27285
rect 20168 27276 20220 27328
rect 23572 27548 23624 27600
rect 24400 27616 24452 27668
rect 26700 27616 26752 27668
rect 27620 27616 27672 27668
rect 25504 27548 25556 27600
rect 28356 27548 28408 27600
rect 22192 27276 22244 27328
rect 23572 27455 23624 27464
rect 23572 27421 23581 27455
rect 23581 27421 23615 27455
rect 23615 27421 23624 27455
rect 23572 27412 23624 27421
rect 29092 27480 29144 27532
rect 29644 27480 29696 27532
rect 28172 27455 28224 27464
rect 28172 27421 28181 27455
rect 28181 27421 28215 27455
rect 28215 27421 28224 27455
rect 28172 27412 28224 27421
rect 26056 27387 26108 27396
rect 26056 27353 26065 27387
rect 26065 27353 26099 27387
rect 26099 27353 26108 27387
rect 26056 27344 26108 27353
rect 27436 27344 27488 27396
rect 29184 27412 29236 27464
rect 30012 27455 30064 27464
rect 30012 27421 30021 27455
rect 30021 27421 30055 27455
rect 30055 27421 30064 27455
rect 30012 27412 30064 27421
rect 30380 27455 30432 27464
rect 30380 27421 30389 27455
rect 30389 27421 30423 27455
rect 30423 27421 30432 27455
rect 30380 27412 30432 27421
rect 30656 27455 30708 27464
rect 30656 27421 30665 27455
rect 30665 27421 30699 27455
rect 30699 27421 30708 27455
rect 30656 27412 30708 27421
rect 30932 27412 30984 27464
rect 34612 27616 34664 27668
rect 33784 27591 33836 27600
rect 33784 27557 33793 27591
rect 33793 27557 33827 27591
rect 33827 27557 33836 27591
rect 33784 27548 33836 27557
rect 34336 27548 34388 27600
rect 26424 27276 26476 27328
rect 27804 27319 27856 27328
rect 27804 27285 27813 27319
rect 27813 27285 27847 27319
rect 27847 27285 27856 27319
rect 27804 27276 27856 27285
rect 27896 27276 27948 27328
rect 28264 27276 28316 27328
rect 32680 27344 32732 27396
rect 29644 27319 29696 27328
rect 29644 27285 29653 27319
rect 29653 27285 29687 27319
rect 29687 27285 29696 27319
rect 29644 27276 29696 27285
rect 29828 27319 29880 27328
rect 29828 27285 29837 27319
rect 29837 27285 29871 27319
rect 29871 27285 29880 27319
rect 29828 27276 29880 27285
rect 30380 27276 30432 27328
rect 31760 27276 31812 27328
rect 33600 27319 33652 27328
rect 33600 27285 33609 27319
rect 33609 27285 33643 27319
rect 33643 27285 33652 27319
rect 33600 27276 33652 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 6828 27072 6880 27124
rect 10048 27072 10100 27124
rect 11612 27072 11664 27124
rect 12164 27072 12216 27124
rect 7196 27004 7248 27056
rect 7380 27004 7432 27056
rect 11888 27004 11940 27056
rect 12256 26979 12308 26988
rect 12256 26945 12265 26979
rect 12265 26945 12299 26979
rect 12299 26945 12308 26979
rect 12256 26936 12308 26945
rect 12348 26979 12400 26988
rect 12348 26945 12358 26979
rect 12358 26945 12392 26979
rect 12392 26945 12400 26979
rect 12348 26936 12400 26945
rect 6920 26911 6972 26920
rect 6920 26877 6929 26911
rect 6929 26877 6963 26911
rect 6963 26877 6972 26911
rect 6920 26868 6972 26877
rect 7472 26868 7524 26920
rect 8392 26911 8444 26920
rect 8392 26877 8401 26911
rect 8401 26877 8435 26911
rect 8435 26877 8444 26911
rect 12808 26936 12860 26988
rect 16304 27072 16356 27124
rect 16672 27115 16724 27124
rect 16672 27081 16681 27115
rect 16681 27081 16715 27115
rect 16715 27081 16724 27115
rect 16672 27072 16724 27081
rect 16948 27115 17000 27124
rect 16948 27081 16957 27115
rect 16957 27081 16991 27115
rect 16991 27081 17000 27115
rect 16948 27072 17000 27081
rect 14004 27004 14056 27056
rect 14372 27004 14424 27056
rect 14648 27004 14700 27056
rect 15476 27047 15528 27056
rect 15476 27013 15485 27047
rect 15485 27013 15519 27047
rect 15519 27013 15528 27047
rect 15476 27004 15528 27013
rect 14740 26979 14792 26988
rect 14740 26945 14749 26979
rect 14749 26945 14783 26979
rect 14783 26945 14792 26979
rect 14740 26936 14792 26945
rect 15016 26936 15068 26988
rect 15384 26936 15436 26988
rect 15660 26979 15712 26988
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 16396 26936 16448 26988
rect 16764 26936 16816 26988
rect 8392 26868 8444 26877
rect 9864 26800 9916 26852
rect 12532 26800 12584 26852
rect 14188 26800 14240 26852
rect 6000 26732 6052 26784
rect 7380 26732 7432 26784
rect 12900 26775 12952 26784
rect 12900 26741 12909 26775
rect 12909 26741 12943 26775
rect 12943 26741 12952 26775
rect 12900 26732 12952 26741
rect 14280 26775 14332 26784
rect 14280 26741 14289 26775
rect 14289 26741 14323 26775
rect 14323 26741 14332 26775
rect 14280 26732 14332 26741
rect 14648 26911 14700 26920
rect 14648 26877 14657 26911
rect 14657 26877 14691 26911
rect 14691 26877 14700 26911
rect 14648 26868 14700 26877
rect 15476 26868 15528 26920
rect 15108 26800 15160 26852
rect 17040 26979 17092 26988
rect 17040 26945 17049 26979
rect 17049 26945 17083 26979
rect 17083 26945 17092 26979
rect 17040 26936 17092 26945
rect 17224 26936 17276 26988
rect 17684 26979 17736 26988
rect 17684 26945 17693 26979
rect 17693 26945 17727 26979
rect 17727 26945 17736 26979
rect 17684 26936 17736 26945
rect 17776 26979 17828 26988
rect 17776 26945 17785 26979
rect 17785 26945 17819 26979
rect 17819 26945 17828 26979
rect 17776 26936 17828 26945
rect 18512 27072 18564 27124
rect 18604 27072 18656 27124
rect 18972 27072 19024 27124
rect 22192 27115 22244 27124
rect 22192 27081 22201 27115
rect 22201 27081 22235 27115
rect 22235 27081 22244 27115
rect 22192 27072 22244 27081
rect 16948 26868 17000 26920
rect 18512 26868 18564 26920
rect 18972 26979 19024 26988
rect 18972 26945 18981 26979
rect 18981 26945 19015 26979
rect 19015 26945 19024 26979
rect 18972 26936 19024 26945
rect 19432 26936 19484 26988
rect 24768 27072 24820 27124
rect 26056 27072 26108 27124
rect 27804 27072 27856 27124
rect 28632 27072 28684 27124
rect 23480 27004 23532 27056
rect 19340 26868 19392 26920
rect 22744 26979 22796 26988
rect 22744 26945 22753 26979
rect 22753 26945 22787 26979
rect 22787 26945 22796 26979
rect 22744 26936 22796 26945
rect 24676 26936 24728 26988
rect 25964 26936 26016 26988
rect 26424 26979 26476 26988
rect 24768 26868 24820 26920
rect 26424 26945 26433 26979
rect 26433 26945 26467 26979
rect 26467 26945 26476 26979
rect 26424 26936 26476 26945
rect 26516 26868 26568 26920
rect 17132 26800 17184 26852
rect 17316 26800 17368 26852
rect 26056 26800 26108 26852
rect 27344 26868 27396 26920
rect 27896 26868 27948 26920
rect 29644 27072 29696 27124
rect 29828 27072 29880 27124
rect 31576 27072 31628 27124
rect 34060 27072 34112 27124
rect 29736 26868 29788 26920
rect 31668 26979 31720 26988
rect 31668 26945 31677 26979
rect 31677 26945 31711 26979
rect 31711 26945 31720 26979
rect 31668 26936 31720 26945
rect 33140 26979 33192 26988
rect 33140 26945 33149 26979
rect 33149 26945 33183 26979
rect 33183 26945 33192 26979
rect 33140 26936 33192 26945
rect 33600 27004 33652 27056
rect 35992 26936 36044 26988
rect 29000 26800 29052 26852
rect 33784 26868 33836 26920
rect 15568 26732 15620 26784
rect 16948 26732 17000 26784
rect 17500 26732 17552 26784
rect 17684 26775 17736 26784
rect 17684 26741 17693 26775
rect 17693 26741 17727 26775
rect 17727 26741 17736 26775
rect 17684 26732 17736 26741
rect 18880 26732 18932 26784
rect 19340 26732 19392 26784
rect 19984 26732 20036 26784
rect 22560 26732 22612 26784
rect 25872 26732 25924 26784
rect 28264 26732 28316 26784
rect 30380 26732 30432 26784
rect 31392 26732 31444 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 6920 26528 6972 26580
rect 12256 26528 12308 26580
rect 13452 26528 13504 26580
rect 14280 26528 14332 26580
rect 14648 26528 14700 26580
rect 7288 26392 7340 26444
rect 11244 26460 11296 26512
rect 7840 26392 7892 26444
rect 8116 26392 8168 26444
rect 8760 26392 8812 26444
rect 14924 26460 14976 26512
rect 5080 26299 5132 26308
rect 5080 26265 5089 26299
rect 5089 26265 5123 26299
rect 5123 26265 5132 26299
rect 5080 26256 5132 26265
rect 3884 26188 3936 26240
rect 6000 26188 6052 26240
rect 6920 26231 6972 26240
rect 6920 26197 6929 26231
rect 6929 26197 6963 26231
rect 6963 26197 6972 26231
rect 6920 26188 6972 26197
rect 7840 26188 7892 26240
rect 8392 26367 8444 26376
rect 8392 26333 8401 26367
rect 8401 26333 8435 26367
rect 8435 26333 8444 26367
rect 8392 26324 8444 26333
rect 12900 26392 12952 26444
rect 8484 26299 8536 26308
rect 8484 26265 8493 26299
rect 8493 26265 8527 26299
rect 8527 26265 8536 26299
rect 8484 26256 8536 26265
rect 8116 26188 8168 26240
rect 9588 26324 9640 26376
rect 11888 26324 11940 26376
rect 12624 26324 12676 26376
rect 14280 26392 14332 26444
rect 13636 26367 13688 26376
rect 13636 26333 13645 26367
rect 13645 26333 13679 26367
rect 13679 26333 13688 26367
rect 13636 26324 13688 26333
rect 14004 26324 14056 26376
rect 17316 26528 17368 26580
rect 17684 26528 17736 26580
rect 18604 26528 18656 26580
rect 19156 26528 19208 26580
rect 15108 26503 15160 26512
rect 15108 26469 15117 26503
rect 15117 26469 15151 26503
rect 15151 26469 15160 26503
rect 15108 26460 15160 26469
rect 15568 26460 15620 26512
rect 14556 26256 14608 26308
rect 15476 26392 15528 26444
rect 15292 26367 15344 26376
rect 15292 26333 15301 26367
rect 15301 26333 15335 26367
rect 15335 26333 15344 26367
rect 15292 26324 15344 26333
rect 15752 26324 15804 26376
rect 16948 26324 17000 26376
rect 8668 26188 8720 26240
rect 12348 26188 12400 26240
rect 15476 26299 15528 26308
rect 15476 26265 15485 26299
rect 15485 26265 15519 26299
rect 15519 26265 15528 26299
rect 15476 26256 15528 26265
rect 15936 26256 15988 26308
rect 17868 26460 17920 26512
rect 17960 26460 18012 26512
rect 22652 26460 22704 26512
rect 17776 26392 17828 26444
rect 25412 26528 25464 26580
rect 25504 26528 25556 26580
rect 17500 26324 17552 26376
rect 20812 26367 20864 26376
rect 20812 26333 20821 26367
rect 20821 26333 20855 26367
rect 20855 26333 20864 26367
rect 20812 26324 20864 26333
rect 20904 26324 20956 26376
rect 17684 26256 17736 26308
rect 20168 26256 20220 26308
rect 20444 26299 20496 26308
rect 20444 26265 20453 26299
rect 20453 26265 20487 26299
rect 20487 26265 20496 26299
rect 20444 26256 20496 26265
rect 22928 26324 22980 26376
rect 23296 26324 23348 26376
rect 24492 26324 24544 26376
rect 21548 26256 21600 26308
rect 24676 26324 24728 26376
rect 25320 26324 25372 26376
rect 25596 26367 25648 26376
rect 25596 26333 25605 26367
rect 25605 26333 25639 26367
rect 25639 26333 25648 26367
rect 25596 26324 25648 26333
rect 26148 26460 26200 26512
rect 28172 26528 28224 26580
rect 30012 26528 30064 26580
rect 33140 26528 33192 26580
rect 26056 26324 26108 26376
rect 26240 26367 26292 26376
rect 26240 26333 26249 26367
rect 26249 26333 26283 26367
rect 26283 26333 26292 26367
rect 26240 26324 26292 26333
rect 26700 26392 26752 26444
rect 29276 26460 29328 26512
rect 28264 26435 28316 26444
rect 28264 26401 28273 26435
rect 28273 26401 28307 26435
rect 28307 26401 28316 26435
rect 28264 26392 28316 26401
rect 28356 26435 28408 26444
rect 28356 26401 28365 26435
rect 28365 26401 28399 26435
rect 28399 26401 28408 26435
rect 28356 26392 28408 26401
rect 30104 26392 30156 26444
rect 29000 26324 29052 26376
rect 30012 26324 30064 26376
rect 30932 26392 30984 26444
rect 31392 26392 31444 26444
rect 32496 26392 32548 26444
rect 33876 26435 33928 26444
rect 33876 26401 33885 26435
rect 33885 26401 33919 26435
rect 33919 26401 33928 26435
rect 33876 26392 33928 26401
rect 30472 26324 30524 26376
rect 32680 26324 32732 26376
rect 33784 26324 33836 26376
rect 34704 26367 34756 26376
rect 34704 26333 34713 26367
rect 34713 26333 34747 26367
rect 34747 26333 34756 26367
rect 34704 26324 34756 26333
rect 34980 26367 35032 26376
rect 34980 26333 34989 26367
rect 34989 26333 35023 26367
rect 35023 26333 35032 26367
rect 34980 26324 35032 26333
rect 29184 26256 29236 26308
rect 31300 26256 31352 26308
rect 31576 26256 31628 26308
rect 32772 26256 32824 26308
rect 34244 26256 34296 26308
rect 35992 26256 36044 26308
rect 36636 26256 36688 26308
rect 17316 26188 17368 26240
rect 20076 26188 20128 26240
rect 22744 26188 22796 26240
rect 23388 26231 23440 26240
rect 23388 26197 23397 26231
rect 23397 26197 23431 26231
rect 23431 26197 23440 26231
rect 23388 26188 23440 26197
rect 23756 26231 23808 26240
rect 23756 26197 23765 26231
rect 23765 26197 23799 26231
rect 23799 26197 23808 26231
rect 23756 26188 23808 26197
rect 26056 26231 26108 26240
rect 26056 26197 26065 26231
rect 26065 26197 26099 26231
rect 26099 26197 26108 26231
rect 26056 26188 26108 26197
rect 27344 26188 27396 26240
rect 27804 26188 27856 26240
rect 32680 26188 32732 26240
rect 33324 26188 33376 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 5080 25984 5132 26036
rect 6920 25984 6972 26036
rect 19248 25984 19300 26036
rect 3884 25916 3936 25968
rect 1768 25891 1820 25900
rect 1768 25857 1777 25891
rect 1777 25857 1811 25891
rect 1811 25857 1820 25891
rect 1768 25848 1820 25857
rect 2964 25848 3016 25900
rect 3056 25891 3108 25900
rect 3056 25857 3065 25891
rect 3065 25857 3099 25891
rect 3099 25857 3108 25891
rect 3056 25848 3108 25857
rect 16764 25916 16816 25968
rect 17776 25916 17828 25968
rect 10048 25848 10100 25900
rect 13820 25848 13872 25900
rect 18420 25916 18472 25968
rect 1860 25780 1912 25832
rect 3608 25823 3660 25832
rect 3608 25789 3617 25823
rect 3617 25789 3651 25823
rect 3651 25789 3660 25823
rect 3608 25780 3660 25789
rect 8668 25823 8720 25832
rect 8668 25789 8677 25823
rect 8677 25789 8711 25823
rect 8711 25789 8720 25823
rect 8668 25780 8720 25789
rect 8944 25823 8996 25832
rect 8944 25789 8953 25823
rect 8953 25789 8987 25823
rect 8987 25789 8996 25823
rect 8944 25780 8996 25789
rect 14648 25780 14700 25832
rect 17960 25848 18012 25900
rect 18328 25848 18380 25900
rect 19800 25984 19852 26036
rect 20812 25984 20864 26036
rect 21180 25984 21232 26036
rect 22468 25984 22520 26036
rect 23756 25984 23808 26036
rect 24768 25984 24820 26036
rect 19892 25916 19944 25968
rect 20260 25916 20312 25968
rect 20536 25916 20588 25968
rect 23020 25916 23072 25968
rect 25136 25984 25188 26036
rect 25320 25984 25372 26036
rect 16580 25780 16632 25832
rect 18144 25780 18196 25832
rect 18420 25780 18472 25832
rect 18972 25848 19024 25900
rect 19340 25891 19392 25900
rect 19340 25857 19358 25891
rect 19358 25857 19392 25891
rect 19340 25848 19392 25857
rect 19800 25891 19852 25900
rect 19800 25857 19809 25891
rect 19809 25857 19843 25891
rect 19843 25857 19852 25891
rect 19800 25848 19852 25857
rect 20444 25891 20496 25900
rect 20444 25857 20453 25891
rect 20453 25857 20487 25891
rect 20487 25857 20496 25891
rect 20444 25848 20496 25857
rect 15108 25712 15160 25764
rect 19524 25712 19576 25764
rect 940 25644 992 25696
rect 2872 25687 2924 25696
rect 2872 25653 2881 25687
rect 2881 25653 2915 25687
rect 2915 25653 2924 25687
rect 2872 25644 2924 25653
rect 5080 25687 5132 25696
rect 5080 25653 5089 25687
rect 5089 25653 5123 25687
rect 5123 25653 5132 25687
rect 5080 25644 5132 25653
rect 9680 25644 9732 25696
rect 13084 25644 13136 25696
rect 18144 25644 18196 25696
rect 19064 25644 19116 25696
rect 19156 25687 19208 25696
rect 19156 25653 19165 25687
rect 19165 25653 19199 25687
rect 19199 25653 19208 25687
rect 19156 25644 19208 25653
rect 19340 25644 19392 25696
rect 20076 25780 20128 25832
rect 19708 25712 19760 25764
rect 20996 25848 21048 25900
rect 22192 25848 22244 25900
rect 22652 25891 22704 25900
rect 22652 25857 22661 25891
rect 22661 25857 22695 25891
rect 22695 25857 22704 25891
rect 22652 25848 22704 25857
rect 20904 25644 20956 25696
rect 20996 25687 21048 25696
rect 20996 25653 21005 25687
rect 21005 25653 21039 25687
rect 21039 25653 21048 25687
rect 20996 25644 21048 25653
rect 21088 25644 21140 25696
rect 21272 25644 21324 25696
rect 22560 25755 22612 25764
rect 22560 25721 22569 25755
rect 22569 25721 22603 25755
rect 22603 25721 22612 25755
rect 22560 25712 22612 25721
rect 22284 25687 22336 25696
rect 22284 25653 22293 25687
rect 22293 25653 22327 25687
rect 22327 25653 22336 25687
rect 22284 25644 22336 25653
rect 22376 25644 22428 25696
rect 23112 25891 23164 25900
rect 23112 25857 23121 25891
rect 23121 25857 23155 25891
rect 23155 25857 23164 25891
rect 23112 25848 23164 25857
rect 22928 25780 22980 25832
rect 23112 25644 23164 25696
rect 23664 25780 23716 25832
rect 24308 25891 24360 25900
rect 24308 25857 24317 25891
rect 24317 25857 24351 25891
rect 24351 25857 24360 25891
rect 24308 25848 24360 25857
rect 24676 25848 24728 25900
rect 24768 25891 24820 25900
rect 24768 25857 24777 25891
rect 24777 25857 24811 25891
rect 24811 25857 24820 25891
rect 24768 25848 24820 25857
rect 23940 25780 23992 25832
rect 24216 25823 24268 25832
rect 24216 25789 24225 25823
rect 24225 25789 24259 25823
rect 24259 25789 24268 25823
rect 24216 25780 24268 25789
rect 25136 25848 25188 25900
rect 25504 25891 25556 25900
rect 25504 25857 25513 25891
rect 25513 25857 25547 25891
rect 25547 25857 25556 25891
rect 25504 25848 25556 25857
rect 26056 25984 26108 26036
rect 29644 25984 29696 26036
rect 30104 25984 30156 26036
rect 31300 25984 31352 26036
rect 25412 25780 25464 25832
rect 24952 25712 25004 25764
rect 25596 25712 25648 25764
rect 31392 25916 31444 25968
rect 31576 26027 31628 26036
rect 31576 25993 31585 26027
rect 31585 25993 31619 26027
rect 31619 25993 31628 26027
rect 31576 25984 31628 25993
rect 31668 25984 31720 26036
rect 32496 25984 32548 26036
rect 34336 25984 34388 26036
rect 34704 25984 34756 26036
rect 34980 25984 35032 26036
rect 26056 25780 26108 25832
rect 26332 25891 26384 25900
rect 26332 25857 26341 25891
rect 26341 25857 26375 25891
rect 26375 25857 26384 25891
rect 26332 25848 26384 25857
rect 27160 25848 27212 25900
rect 31760 25891 31812 25900
rect 31760 25857 31769 25891
rect 31769 25857 31803 25891
rect 31803 25857 31812 25891
rect 31760 25848 31812 25857
rect 32772 25848 32824 25900
rect 28632 25780 28684 25832
rect 30656 25780 30708 25832
rect 32680 25823 32732 25832
rect 32680 25789 32689 25823
rect 32689 25789 32723 25823
rect 32723 25789 32732 25823
rect 32680 25780 32732 25789
rect 25964 25712 26016 25764
rect 26332 25712 26384 25764
rect 24124 25687 24176 25696
rect 24124 25653 24133 25687
rect 24133 25653 24167 25687
rect 24167 25653 24176 25687
rect 24124 25644 24176 25653
rect 25320 25687 25372 25696
rect 25320 25653 25329 25687
rect 25329 25653 25363 25687
rect 25363 25653 25372 25687
rect 25320 25644 25372 25653
rect 26608 25687 26660 25696
rect 26608 25653 26617 25687
rect 26617 25653 26651 25687
rect 26651 25653 26660 25687
rect 26608 25644 26660 25653
rect 27528 25644 27580 25696
rect 30012 25644 30064 25696
rect 30288 25644 30340 25696
rect 33232 25891 33284 25900
rect 33232 25857 33241 25891
rect 33241 25857 33275 25891
rect 33275 25857 33284 25891
rect 33232 25848 33284 25857
rect 33324 25891 33376 25900
rect 33324 25857 33333 25891
rect 33333 25857 33367 25891
rect 33367 25857 33376 25891
rect 33324 25848 33376 25857
rect 34152 25823 34204 25832
rect 34152 25789 34161 25823
rect 34161 25789 34195 25823
rect 34195 25789 34204 25823
rect 34152 25780 34204 25789
rect 34244 25780 34296 25832
rect 36636 25848 36688 25900
rect 34704 25712 34756 25764
rect 34796 25644 34848 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3608 25440 3660 25492
rect 8944 25440 8996 25492
rect 9680 25440 9732 25492
rect 2872 25304 2924 25356
rect 1400 25236 1452 25288
rect 1860 25279 1912 25288
rect 1860 25245 1869 25279
rect 1869 25245 1903 25279
rect 1903 25245 1912 25279
rect 1860 25236 1912 25245
rect 4344 25236 4396 25288
rect 7564 25279 7616 25288
rect 7564 25245 7573 25279
rect 7573 25245 7607 25279
rect 7607 25245 7616 25279
rect 7564 25236 7616 25245
rect 9864 25347 9916 25356
rect 9864 25313 9873 25347
rect 9873 25313 9907 25347
rect 9907 25313 9916 25347
rect 9864 25304 9916 25313
rect 2872 25168 2924 25220
rect 9036 25168 9088 25220
rect 4620 25100 4672 25152
rect 7288 25100 7340 25152
rect 10140 25279 10192 25288
rect 10140 25245 10149 25279
rect 10149 25245 10183 25279
rect 10183 25245 10192 25279
rect 10140 25236 10192 25245
rect 13084 25440 13136 25492
rect 19248 25440 19300 25492
rect 20444 25440 20496 25492
rect 12256 25304 12308 25356
rect 13176 25304 13228 25356
rect 12624 25236 12676 25288
rect 13084 25279 13136 25288
rect 13084 25245 13093 25279
rect 13093 25245 13127 25279
rect 13127 25245 13136 25279
rect 13084 25236 13136 25245
rect 15108 25372 15160 25424
rect 15200 25372 15252 25424
rect 17132 25372 17184 25424
rect 14832 25347 14884 25356
rect 14832 25313 14841 25347
rect 14841 25313 14875 25347
rect 14875 25313 14884 25347
rect 14832 25304 14884 25313
rect 13452 25279 13504 25288
rect 13452 25245 13461 25279
rect 13461 25245 13495 25279
rect 13495 25245 13504 25279
rect 13452 25236 13504 25245
rect 10508 25168 10560 25220
rect 11060 25168 11112 25220
rect 11796 25168 11848 25220
rect 12532 25168 12584 25220
rect 14188 25168 14240 25220
rect 15660 25236 15712 25288
rect 16212 25236 16264 25288
rect 9588 25100 9640 25152
rect 11980 25143 12032 25152
rect 11980 25109 11989 25143
rect 11989 25109 12023 25143
rect 12023 25109 12032 25143
rect 11980 25100 12032 25109
rect 12348 25100 12400 25152
rect 12808 25100 12860 25152
rect 16948 25236 17000 25288
rect 17040 25279 17092 25288
rect 17040 25245 17049 25279
rect 17049 25245 17083 25279
rect 17083 25245 17092 25279
rect 17040 25236 17092 25245
rect 17868 25372 17920 25424
rect 22468 25440 22520 25492
rect 22560 25440 22612 25492
rect 23572 25440 23624 25492
rect 24768 25483 24820 25492
rect 24768 25449 24777 25483
rect 24777 25449 24811 25483
rect 24811 25449 24820 25483
rect 24768 25440 24820 25449
rect 18144 25304 18196 25356
rect 20904 25372 20956 25424
rect 20996 25347 21048 25356
rect 20996 25313 21005 25347
rect 21005 25313 21039 25347
rect 21039 25313 21048 25347
rect 20996 25304 21048 25313
rect 18236 25236 18288 25288
rect 18512 25279 18564 25288
rect 18512 25245 18521 25279
rect 18521 25245 18555 25279
rect 18555 25245 18564 25279
rect 18512 25236 18564 25245
rect 20720 25279 20772 25288
rect 20720 25245 20729 25279
rect 20729 25245 20763 25279
rect 20763 25245 20772 25279
rect 20720 25236 20772 25245
rect 20076 25168 20128 25220
rect 20352 25168 20404 25220
rect 16764 25100 16816 25152
rect 17132 25100 17184 25152
rect 17868 25100 17920 25152
rect 19892 25100 19944 25152
rect 20628 25100 20680 25152
rect 21272 25372 21324 25424
rect 21180 25236 21232 25288
rect 21456 25279 21508 25288
rect 21456 25245 21465 25279
rect 21465 25245 21499 25279
rect 21499 25245 21508 25279
rect 21456 25236 21508 25245
rect 21732 25279 21784 25288
rect 21732 25245 21741 25279
rect 21741 25245 21775 25279
rect 21775 25245 21784 25279
rect 21732 25236 21784 25245
rect 21180 25100 21232 25152
rect 22008 25168 22060 25220
rect 22192 25279 22244 25288
rect 22192 25245 22201 25279
rect 22201 25245 22235 25279
rect 22235 25245 22244 25279
rect 22192 25236 22244 25245
rect 22376 25279 22428 25288
rect 22376 25245 22383 25279
rect 22383 25245 22428 25279
rect 22376 25236 22428 25245
rect 22652 25372 22704 25424
rect 24216 25372 24268 25424
rect 26884 25440 26936 25492
rect 31852 25440 31904 25492
rect 33324 25440 33376 25492
rect 23112 25304 23164 25356
rect 23480 25347 23532 25356
rect 23480 25313 23489 25347
rect 23489 25313 23523 25347
rect 23523 25313 23532 25347
rect 23480 25304 23532 25313
rect 26240 25372 26292 25424
rect 26424 25372 26476 25424
rect 26148 25304 26200 25356
rect 22468 25211 22520 25220
rect 22468 25177 22477 25211
rect 22477 25177 22511 25211
rect 22511 25177 22520 25211
rect 22468 25168 22520 25177
rect 22652 25100 22704 25152
rect 22744 25100 22796 25152
rect 25320 25100 25372 25152
rect 26056 25236 26108 25288
rect 26792 25236 26844 25288
rect 27528 25304 27580 25356
rect 27896 25372 27948 25424
rect 28908 25372 28960 25424
rect 27528 25211 27580 25220
rect 27528 25177 27537 25211
rect 27537 25177 27571 25211
rect 27571 25177 27580 25211
rect 27528 25168 27580 25177
rect 26700 25100 26752 25152
rect 27160 25100 27212 25152
rect 28264 25236 28316 25288
rect 28632 25236 28684 25288
rect 29092 25304 29144 25356
rect 34704 25372 34756 25424
rect 30104 25168 30156 25220
rect 30932 25236 30984 25288
rect 34336 25279 34388 25288
rect 34336 25245 34345 25279
rect 34345 25245 34379 25279
rect 34379 25245 34388 25279
rect 34336 25236 34388 25245
rect 29092 25143 29144 25152
rect 29092 25109 29101 25143
rect 29101 25109 29135 25143
rect 29135 25109 29144 25143
rect 29092 25100 29144 25109
rect 30288 25100 30340 25152
rect 31300 25100 31352 25152
rect 35992 25168 36044 25220
rect 36728 25211 36780 25220
rect 36728 25177 36737 25211
rect 36737 25177 36771 25211
rect 36771 25177 36780 25211
rect 36728 25168 36780 25177
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4344 24939 4396 24948
rect 4344 24905 4353 24939
rect 4353 24905 4387 24939
rect 4387 24905 4396 24939
rect 4344 24896 4396 24905
rect 5080 24896 5132 24948
rect 5816 24896 5868 24948
rect 9220 24939 9272 24948
rect 9220 24905 9229 24939
rect 9229 24905 9263 24939
rect 9263 24905 9272 24939
rect 9220 24896 9272 24905
rect 9588 24939 9640 24948
rect 9588 24905 9597 24939
rect 9597 24905 9631 24939
rect 9631 24905 9640 24939
rect 9588 24896 9640 24905
rect 10140 24896 10192 24948
rect 10508 24896 10560 24948
rect 11980 24896 12032 24948
rect 6000 24828 6052 24880
rect 5908 24803 5960 24812
rect 5908 24769 5917 24803
rect 5917 24769 5951 24803
rect 5951 24769 5960 24803
rect 5908 24760 5960 24769
rect 10416 24803 10468 24812
rect 10416 24769 10425 24803
rect 10425 24769 10459 24803
rect 10459 24769 10468 24803
rect 10416 24760 10468 24769
rect 12348 24871 12400 24880
rect 12348 24837 12357 24871
rect 12357 24837 12391 24871
rect 12391 24837 12400 24871
rect 12348 24828 12400 24837
rect 14188 24896 14240 24948
rect 13176 24828 13228 24880
rect 15200 24896 15252 24948
rect 16948 24896 17000 24948
rect 12256 24760 12308 24812
rect 1400 24735 1452 24744
rect 1400 24701 1409 24735
rect 1409 24701 1443 24735
rect 1443 24701 1452 24735
rect 1400 24692 1452 24701
rect 1676 24735 1728 24744
rect 1676 24701 1685 24735
rect 1685 24701 1719 24735
rect 1719 24701 1728 24735
rect 1676 24692 1728 24701
rect 2872 24692 2924 24744
rect 4804 24735 4856 24744
rect 4804 24701 4813 24735
rect 4813 24701 4847 24735
rect 4847 24701 4856 24735
rect 4804 24692 4856 24701
rect 3148 24599 3200 24608
rect 3148 24565 3157 24599
rect 3157 24565 3191 24599
rect 3191 24565 3200 24599
rect 3148 24556 3200 24565
rect 3976 24556 4028 24608
rect 7288 24735 7340 24744
rect 7288 24701 7297 24735
rect 7297 24701 7331 24735
rect 7331 24701 7340 24735
rect 7288 24692 7340 24701
rect 7932 24692 7984 24744
rect 9864 24735 9916 24744
rect 9864 24701 9873 24735
rect 9873 24701 9907 24735
rect 9907 24701 9916 24735
rect 9864 24692 9916 24701
rect 13544 24760 13596 24812
rect 14556 24828 14608 24880
rect 15752 24828 15804 24880
rect 16304 24828 16356 24880
rect 5632 24556 5684 24608
rect 7104 24556 7156 24608
rect 12532 24556 12584 24608
rect 14556 24692 14608 24744
rect 14740 24692 14792 24744
rect 15384 24803 15436 24812
rect 15384 24769 15393 24803
rect 15393 24769 15427 24803
rect 15427 24769 15436 24803
rect 15384 24760 15436 24769
rect 16764 24828 16816 24880
rect 17592 24896 17644 24948
rect 17132 24760 17184 24812
rect 17684 24828 17736 24880
rect 18236 24828 18288 24880
rect 18604 24896 18656 24948
rect 18880 24896 18932 24948
rect 22928 24896 22980 24948
rect 23020 24896 23072 24948
rect 27528 24896 27580 24948
rect 29092 24896 29144 24948
rect 30104 24896 30156 24948
rect 20996 24828 21048 24880
rect 21088 24871 21140 24880
rect 21088 24837 21097 24871
rect 21097 24837 21131 24871
rect 21131 24837 21140 24871
rect 21088 24828 21140 24837
rect 14924 24692 14976 24744
rect 13176 24599 13228 24608
rect 13176 24565 13185 24599
rect 13185 24565 13219 24599
rect 13219 24565 13228 24599
rect 13176 24556 13228 24565
rect 14096 24556 14148 24608
rect 15108 24556 15160 24608
rect 16856 24624 16908 24676
rect 19800 24760 19852 24812
rect 20076 24760 20128 24812
rect 22008 24828 22060 24880
rect 25412 24828 25464 24880
rect 26424 24828 26476 24880
rect 27344 24871 27396 24880
rect 27344 24837 27353 24871
rect 27353 24837 27387 24871
rect 27387 24837 27396 24871
rect 27344 24828 27396 24837
rect 21548 24760 21600 24812
rect 21732 24760 21784 24812
rect 22652 24760 22704 24812
rect 23480 24803 23532 24812
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 23572 24760 23624 24812
rect 25136 24760 25188 24812
rect 25872 24803 25924 24812
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 17684 24692 17736 24744
rect 17868 24735 17920 24744
rect 17868 24701 17877 24735
rect 17877 24701 17911 24735
rect 17911 24701 17920 24735
rect 17868 24692 17920 24701
rect 20444 24692 20496 24744
rect 22192 24692 22244 24744
rect 23848 24692 23900 24744
rect 25412 24692 25464 24744
rect 17408 24624 17460 24676
rect 17960 24624 18012 24676
rect 19340 24624 19392 24676
rect 24216 24624 24268 24676
rect 28816 24760 28868 24812
rect 29644 24828 29696 24880
rect 30932 24871 30984 24880
rect 30932 24837 30941 24871
rect 30941 24837 30975 24871
rect 30975 24837 30984 24871
rect 30932 24828 30984 24837
rect 31116 24803 31168 24812
rect 31116 24769 31125 24803
rect 31125 24769 31159 24803
rect 31159 24769 31168 24803
rect 31116 24760 31168 24769
rect 33232 24896 33284 24948
rect 33324 24896 33376 24948
rect 34336 24896 34388 24948
rect 31852 24828 31904 24880
rect 36728 24828 36780 24880
rect 18512 24599 18564 24608
rect 18512 24565 18521 24599
rect 18521 24565 18555 24599
rect 18555 24565 18564 24599
rect 18512 24556 18564 24565
rect 19524 24556 19576 24608
rect 21272 24556 21324 24608
rect 21364 24556 21416 24608
rect 25504 24556 25556 24608
rect 25964 24599 26016 24608
rect 25964 24565 25973 24599
rect 25973 24565 26007 24599
rect 26007 24565 26016 24599
rect 25964 24556 26016 24565
rect 27804 24692 27856 24744
rect 29736 24692 29788 24744
rect 33048 24692 33100 24744
rect 33140 24692 33192 24744
rect 33784 24760 33836 24812
rect 33324 24692 33376 24744
rect 30288 24624 30340 24676
rect 29000 24556 29052 24608
rect 30196 24556 30248 24608
rect 31208 24599 31260 24608
rect 31208 24565 31217 24599
rect 31217 24565 31251 24599
rect 31251 24565 31260 24599
rect 31208 24556 31260 24565
rect 33324 24556 33376 24608
rect 33416 24556 33468 24608
rect 34152 24556 34204 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1676 24352 1728 24404
rect 3056 24352 3108 24404
rect 4068 24352 4120 24404
rect 7840 24352 7892 24404
rect 7932 24395 7984 24404
rect 7932 24361 7941 24395
rect 7941 24361 7975 24395
rect 7975 24361 7984 24395
rect 7932 24352 7984 24361
rect 9220 24352 9272 24404
rect 1400 24284 1452 24336
rect 3240 24216 3292 24268
rect 3976 24216 4028 24268
rect 5632 24216 5684 24268
rect 15384 24352 15436 24404
rect 15844 24352 15896 24404
rect 14740 24284 14792 24336
rect 15200 24327 15252 24336
rect 15200 24293 15209 24327
rect 15209 24293 15243 24327
rect 15243 24293 15252 24327
rect 15200 24284 15252 24293
rect 15568 24284 15620 24336
rect 4620 24148 4672 24200
rect 12716 24216 12768 24268
rect 13728 24216 13780 24268
rect 9128 24191 9180 24200
rect 9128 24157 9137 24191
rect 9137 24157 9171 24191
rect 9171 24157 9180 24191
rect 9128 24148 9180 24157
rect 3148 24080 3200 24132
rect 6000 24080 6052 24132
rect 15292 24216 15344 24268
rect 16764 24216 16816 24268
rect 18328 24352 18380 24404
rect 19156 24352 19208 24404
rect 17132 24284 17184 24336
rect 17316 24284 17368 24336
rect 17960 24284 18012 24336
rect 18696 24284 18748 24336
rect 23664 24352 23716 24404
rect 25412 24352 25464 24404
rect 25504 24352 25556 24404
rect 14924 24148 14976 24200
rect 15108 24148 15160 24200
rect 14556 24080 14608 24132
rect 15016 24080 15068 24132
rect 15844 24148 15896 24200
rect 16028 24191 16080 24200
rect 16028 24157 16037 24191
rect 16037 24157 16071 24191
rect 16071 24157 16080 24191
rect 16028 24148 16080 24157
rect 16948 24080 17000 24132
rect 17500 24191 17552 24200
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 17500 24148 17552 24157
rect 17868 24191 17920 24200
rect 17868 24157 17877 24191
rect 17877 24157 17911 24191
rect 17911 24157 17920 24191
rect 17868 24148 17920 24157
rect 18236 24148 18288 24200
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 17408 24080 17460 24132
rect 20352 24284 20404 24336
rect 22100 24327 22152 24336
rect 22100 24293 22109 24327
rect 22109 24293 22143 24327
rect 22143 24293 22152 24327
rect 22100 24284 22152 24293
rect 19156 24216 19208 24268
rect 19064 24191 19116 24200
rect 19064 24157 19073 24191
rect 19073 24157 19107 24191
rect 19107 24157 19116 24191
rect 19064 24148 19116 24157
rect 19432 24148 19484 24200
rect 19800 24216 19852 24268
rect 19984 24191 20036 24200
rect 19984 24157 19993 24191
rect 19993 24157 20027 24191
rect 20027 24157 20036 24191
rect 22008 24216 22060 24268
rect 22652 24216 22704 24268
rect 23572 24284 23624 24336
rect 24676 24284 24728 24336
rect 26976 24284 27028 24336
rect 27528 24352 27580 24404
rect 31208 24352 31260 24404
rect 19984 24148 20036 24157
rect 2780 24055 2832 24064
rect 2780 24021 2789 24055
rect 2789 24021 2823 24055
rect 2823 24021 2832 24055
rect 2780 24012 2832 24021
rect 4620 24012 4672 24064
rect 6920 24012 6972 24064
rect 9036 24055 9088 24064
rect 9036 24021 9045 24055
rect 9045 24021 9079 24055
rect 9079 24021 9088 24055
rect 9036 24012 9088 24021
rect 12624 24055 12676 24064
rect 12624 24021 12633 24055
rect 12633 24021 12667 24055
rect 12667 24021 12676 24055
rect 12624 24012 12676 24021
rect 13912 24012 13964 24064
rect 15476 24012 15528 24064
rect 19156 24080 19208 24132
rect 20444 24191 20496 24200
rect 20444 24157 20453 24191
rect 20453 24157 20487 24191
rect 20487 24157 20496 24191
rect 20444 24148 20496 24157
rect 20536 24191 20588 24200
rect 20536 24157 20545 24191
rect 20545 24157 20579 24191
rect 20579 24157 20588 24191
rect 20536 24148 20588 24157
rect 23480 24148 23532 24200
rect 23756 24148 23808 24200
rect 23940 24191 23992 24200
rect 23940 24157 23949 24191
rect 23949 24157 23983 24191
rect 23983 24157 23992 24191
rect 23940 24148 23992 24157
rect 24216 24191 24268 24200
rect 24216 24157 24225 24191
rect 24225 24157 24259 24191
rect 24259 24157 24268 24191
rect 24216 24148 24268 24157
rect 25964 24216 26016 24268
rect 27344 24216 27396 24268
rect 25320 24191 25372 24200
rect 25320 24157 25329 24191
rect 25329 24157 25363 24191
rect 25363 24157 25372 24191
rect 25320 24148 25372 24157
rect 28172 24191 28224 24200
rect 28172 24157 28181 24191
rect 28181 24157 28215 24191
rect 28215 24157 28224 24191
rect 28172 24148 28224 24157
rect 28448 24191 28500 24200
rect 28448 24157 28457 24191
rect 28457 24157 28491 24191
rect 28491 24157 28500 24191
rect 28448 24148 28500 24157
rect 29460 24148 29512 24200
rect 29736 24191 29788 24200
rect 29736 24157 29740 24191
rect 29740 24157 29774 24191
rect 29774 24157 29788 24191
rect 29736 24148 29788 24157
rect 30104 24284 30156 24336
rect 29920 24191 29972 24200
rect 29920 24157 29929 24191
rect 29929 24157 29963 24191
rect 29963 24157 29972 24191
rect 29920 24148 29972 24157
rect 33508 24327 33560 24336
rect 33508 24293 33517 24327
rect 33517 24293 33551 24327
rect 33551 24293 33560 24327
rect 33508 24284 33560 24293
rect 33048 24259 33100 24268
rect 33048 24225 33057 24259
rect 33057 24225 33091 24259
rect 33091 24225 33100 24259
rect 33048 24216 33100 24225
rect 27436 24080 27488 24132
rect 32772 24191 32824 24200
rect 32772 24157 32781 24191
rect 32781 24157 32815 24191
rect 32815 24157 32824 24191
rect 32772 24148 32824 24157
rect 32956 24148 33008 24200
rect 33140 24191 33192 24200
rect 33140 24157 33149 24191
rect 33149 24157 33183 24191
rect 33183 24157 33192 24191
rect 33140 24148 33192 24157
rect 33324 24191 33376 24200
rect 33324 24157 33333 24191
rect 33333 24157 33367 24191
rect 33367 24157 33376 24191
rect 33324 24148 33376 24157
rect 33784 24148 33836 24200
rect 19064 24012 19116 24064
rect 19248 24055 19300 24064
rect 19248 24021 19257 24055
rect 19257 24021 19291 24055
rect 19291 24021 19300 24055
rect 19248 24012 19300 24021
rect 20168 24012 20220 24064
rect 22192 24012 22244 24064
rect 26516 24012 26568 24064
rect 27620 24012 27672 24064
rect 30196 24055 30248 24064
rect 30196 24021 30205 24055
rect 30205 24021 30239 24055
rect 30239 24021 30248 24055
rect 30196 24012 30248 24021
rect 31484 24055 31536 24064
rect 31484 24021 31493 24055
rect 31493 24021 31527 24055
rect 31527 24021 31536 24055
rect 31484 24012 31536 24021
rect 32404 24055 32456 24064
rect 32404 24021 32413 24055
rect 32413 24021 32447 24055
rect 32447 24021 32456 24055
rect 32404 24012 32456 24021
rect 32588 24055 32640 24064
rect 32588 24021 32597 24055
rect 32597 24021 32631 24055
rect 32631 24021 32640 24055
rect 32588 24012 32640 24021
rect 33140 24012 33192 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1952 23808 2004 23860
rect 5908 23808 5960 23860
rect 6920 23808 6972 23860
rect 7288 23808 7340 23860
rect 5632 23715 5684 23724
rect 5632 23681 5641 23715
rect 5641 23681 5675 23715
rect 5675 23681 5684 23715
rect 5632 23672 5684 23681
rect 7012 23672 7064 23724
rect 3976 23604 4028 23656
rect 6000 23536 6052 23588
rect 7288 23536 7340 23588
rect 5264 23468 5316 23520
rect 9036 23740 9088 23792
rect 9956 23808 10008 23860
rect 14832 23808 14884 23860
rect 15660 23808 15712 23860
rect 15936 23808 15988 23860
rect 16948 23808 17000 23860
rect 17040 23808 17092 23860
rect 12716 23740 12768 23792
rect 13452 23783 13504 23792
rect 13452 23749 13461 23783
rect 13461 23749 13495 23783
rect 13495 23749 13504 23783
rect 13452 23740 13504 23749
rect 13912 23740 13964 23792
rect 14280 23783 14332 23792
rect 14280 23749 14289 23783
rect 14289 23749 14323 23783
rect 14323 23749 14332 23783
rect 14280 23740 14332 23749
rect 14464 23740 14516 23792
rect 15016 23783 15068 23792
rect 15016 23749 15025 23783
rect 15025 23749 15059 23783
rect 15059 23749 15068 23783
rect 15016 23740 15068 23749
rect 11152 23715 11204 23724
rect 11152 23681 11161 23715
rect 11161 23681 11195 23715
rect 11195 23681 11204 23715
rect 11152 23672 11204 23681
rect 12900 23715 12952 23724
rect 12900 23681 12909 23715
rect 12909 23681 12943 23715
rect 12943 23681 12952 23715
rect 12900 23672 12952 23681
rect 12992 23715 13044 23724
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 14188 23715 14240 23724
rect 14188 23681 14197 23715
rect 14197 23681 14231 23715
rect 14231 23681 14240 23715
rect 14188 23672 14240 23681
rect 9312 23604 9364 23656
rect 10048 23536 10100 23588
rect 12532 23604 12584 23656
rect 13728 23604 13780 23656
rect 14924 23672 14976 23724
rect 15108 23672 15160 23724
rect 15292 23715 15344 23724
rect 15292 23681 15301 23715
rect 15301 23681 15335 23715
rect 15335 23681 15344 23715
rect 15292 23672 15344 23681
rect 15476 23715 15528 23724
rect 15476 23681 15485 23715
rect 15485 23681 15519 23715
rect 15519 23681 15528 23715
rect 15476 23672 15528 23681
rect 14556 23604 14608 23656
rect 16856 23740 16908 23792
rect 16764 23672 16816 23724
rect 17776 23740 17828 23792
rect 17684 23672 17736 23724
rect 16028 23604 16080 23656
rect 17500 23647 17552 23656
rect 17500 23613 17509 23647
rect 17509 23613 17543 23647
rect 17543 23613 17552 23647
rect 18696 23851 18748 23860
rect 18696 23817 18705 23851
rect 18705 23817 18739 23851
rect 18739 23817 18748 23851
rect 18696 23808 18748 23817
rect 19248 23808 19300 23860
rect 19340 23851 19392 23860
rect 19340 23817 19349 23851
rect 19349 23817 19383 23851
rect 19383 23817 19392 23851
rect 19340 23808 19392 23817
rect 19708 23808 19760 23860
rect 20536 23808 20588 23860
rect 23112 23808 23164 23860
rect 23388 23808 23440 23860
rect 19156 23715 19208 23724
rect 19156 23681 19165 23715
rect 19165 23681 19199 23715
rect 19199 23681 19208 23715
rect 19156 23672 19208 23681
rect 19340 23672 19392 23724
rect 19524 23672 19576 23724
rect 20168 23740 20220 23792
rect 20260 23740 20312 23792
rect 17500 23604 17552 23613
rect 14832 23468 14884 23520
rect 16212 23468 16264 23520
rect 17316 23536 17368 23588
rect 17592 23468 17644 23520
rect 17776 23511 17828 23520
rect 17776 23477 17785 23511
rect 17785 23477 17819 23511
rect 17819 23477 17828 23511
rect 17776 23468 17828 23477
rect 18420 23536 18472 23588
rect 19892 23536 19944 23588
rect 21364 23740 21416 23792
rect 22652 23740 22704 23792
rect 20812 23715 20864 23724
rect 20812 23681 20821 23715
rect 20821 23681 20855 23715
rect 20855 23681 20864 23715
rect 20812 23672 20864 23681
rect 22928 23672 22980 23724
rect 23020 23672 23072 23724
rect 23756 23672 23808 23724
rect 23848 23715 23900 23724
rect 23848 23681 23857 23715
rect 23857 23681 23891 23715
rect 23891 23681 23900 23715
rect 23848 23672 23900 23681
rect 25320 23740 25372 23792
rect 24768 23672 24820 23724
rect 25136 23715 25188 23724
rect 25136 23681 25145 23715
rect 25145 23681 25179 23715
rect 25179 23681 25188 23715
rect 25136 23672 25188 23681
rect 26056 23715 26108 23724
rect 26056 23681 26065 23715
rect 26065 23681 26099 23715
rect 26099 23681 26108 23715
rect 26056 23672 26108 23681
rect 26424 23808 26476 23860
rect 28816 23808 28868 23860
rect 31484 23808 31536 23860
rect 20352 23536 20404 23588
rect 22192 23579 22244 23588
rect 22192 23545 22201 23579
rect 22201 23545 22235 23579
rect 22235 23545 22244 23579
rect 24400 23604 24452 23656
rect 25872 23604 25924 23656
rect 27160 23740 27212 23792
rect 27068 23715 27120 23724
rect 27068 23681 27077 23715
rect 27077 23681 27111 23715
rect 27111 23681 27120 23715
rect 27068 23672 27120 23681
rect 27528 23672 27580 23724
rect 27712 23715 27764 23724
rect 27712 23681 27721 23715
rect 27721 23681 27755 23715
rect 27755 23681 27764 23715
rect 27712 23672 27764 23681
rect 28172 23740 28224 23792
rect 28908 23740 28960 23792
rect 32956 23808 33008 23860
rect 33140 23808 33192 23860
rect 22192 23536 22244 23545
rect 24308 23579 24360 23588
rect 24308 23545 24317 23579
rect 24317 23545 24351 23579
rect 24351 23545 24360 23579
rect 24308 23536 24360 23545
rect 19800 23468 19852 23520
rect 27160 23536 27212 23588
rect 27436 23536 27488 23588
rect 27620 23579 27672 23588
rect 27620 23545 27629 23579
rect 27629 23545 27663 23579
rect 27663 23545 27672 23579
rect 27620 23536 27672 23545
rect 27712 23536 27764 23588
rect 34612 23672 34664 23724
rect 33416 23604 33468 23656
rect 35348 23604 35400 23656
rect 35808 23647 35860 23656
rect 35808 23613 35817 23647
rect 35817 23613 35851 23647
rect 35851 23613 35860 23647
rect 35808 23604 35860 23613
rect 33048 23536 33100 23588
rect 33232 23511 33284 23520
rect 33232 23477 33241 23511
rect 33241 23477 33275 23511
rect 33275 23477 33284 23511
rect 33232 23468 33284 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1768 23264 1820 23316
rect 2780 23264 2832 23316
rect 1952 23103 2004 23112
rect 1952 23069 1961 23103
rect 1961 23069 1995 23103
rect 1995 23069 2004 23103
rect 1952 23060 2004 23069
rect 2688 23103 2740 23112
rect 2688 23069 2697 23103
rect 2697 23069 2731 23103
rect 2731 23069 2740 23103
rect 2688 23060 2740 23069
rect 4160 23264 4212 23316
rect 4620 23264 4672 23316
rect 4804 23264 4856 23316
rect 5632 23264 5684 23316
rect 3148 23103 3200 23112
rect 3148 23069 3157 23103
rect 3157 23069 3191 23103
rect 3191 23069 3200 23103
rect 3148 23060 3200 23069
rect 3608 23103 3660 23112
rect 3608 23069 3617 23103
rect 3617 23069 3651 23103
rect 3651 23069 3660 23103
rect 3608 23060 3660 23069
rect 4436 23103 4488 23112
rect 4436 23069 4445 23103
rect 4445 23069 4479 23103
rect 4479 23069 4488 23103
rect 4436 23060 4488 23069
rect 5356 23196 5408 23248
rect 5816 23196 5868 23248
rect 7012 23307 7064 23316
rect 7012 23273 7021 23307
rect 7021 23273 7055 23307
rect 7055 23273 7064 23307
rect 7012 23264 7064 23273
rect 7196 23264 7248 23316
rect 9312 23307 9364 23316
rect 9312 23273 9321 23307
rect 9321 23273 9355 23307
rect 9355 23273 9364 23307
rect 9312 23264 9364 23273
rect 9404 23264 9456 23316
rect 4896 23103 4948 23112
rect 4896 23069 4905 23103
rect 4905 23069 4939 23103
rect 4939 23069 4948 23103
rect 4896 23060 4948 23069
rect 6552 23128 6604 23180
rect 5908 23103 5960 23112
rect 5908 23069 5917 23103
rect 5917 23069 5951 23103
rect 5951 23069 5960 23103
rect 5908 23060 5960 23069
rect 10140 23196 10192 23248
rect 10600 23196 10652 23248
rect 14188 23264 14240 23316
rect 15016 23264 15068 23316
rect 15292 23264 15344 23316
rect 16028 23264 16080 23316
rect 19800 23264 19852 23316
rect 19892 23264 19944 23316
rect 20812 23307 20864 23316
rect 20812 23273 20821 23307
rect 20821 23273 20855 23307
rect 20855 23273 20864 23307
rect 20812 23264 20864 23273
rect 1860 22924 1912 22976
rect 2504 22924 2556 22976
rect 2872 22924 2924 22976
rect 3976 22924 4028 22976
rect 4528 23035 4580 23044
rect 4528 23001 4537 23035
rect 4537 23001 4571 23035
rect 4571 23001 4580 23035
rect 4528 22992 4580 23001
rect 5264 23035 5316 23044
rect 5264 23001 5273 23035
rect 5273 23001 5307 23035
rect 5307 23001 5316 23035
rect 5264 22992 5316 23001
rect 5356 23035 5408 23044
rect 5356 23001 5365 23035
rect 5365 23001 5399 23035
rect 5399 23001 5408 23035
rect 5356 22992 5408 23001
rect 4620 22924 4672 22976
rect 7012 23060 7064 23112
rect 9128 23128 9180 23180
rect 6000 22924 6052 22976
rect 7196 22992 7248 23044
rect 7380 23035 7432 23044
rect 7380 23001 7389 23035
rect 7389 23001 7423 23035
rect 7423 23001 7432 23035
rect 7380 22992 7432 23001
rect 7564 22992 7616 23044
rect 9404 23060 9456 23112
rect 9496 23103 9548 23112
rect 9496 23069 9505 23103
rect 9505 23069 9539 23103
rect 9539 23069 9548 23103
rect 9496 23060 9548 23069
rect 7932 23035 7984 23044
rect 7932 23001 7941 23035
rect 7941 23001 7975 23035
rect 7975 23001 7984 23035
rect 7932 22992 7984 23001
rect 9680 23035 9732 23044
rect 9680 23001 9689 23035
rect 9689 23001 9723 23035
rect 9723 23001 9732 23035
rect 9680 22992 9732 23001
rect 9864 23103 9916 23112
rect 9864 23069 9873 23103
rect 9873 23069 9907 23103
rect 9907 23069 9916 23103
rect 9864 23060 9916 23069
rect 10048 23060 10100 23112
rect 11152 23128 11204 23180
rect 12072 23128 12124 23180
rect 12348 23128 12400 23180
rect 15568 23128 15620 23180
rect 15660 23171 15712 23180
rect 15660 23137 15669 23171
rect 15669 23137 15703 23171
rect 15703 23137 15712 23171
rect 15660 23128 15712 23137
rect 16120 23128 16172 23180
rect 12716 23060 12768 23112
rect 15016 23060 15068 23112
rect 15108 23060 15160 23112
rect 15384 23103 15436 23112
rect 15384 23069 15393 23103
rect 15393 23069 15427 23103
rect 15427 23069 15436 23103
rect 15384 23060 15436 23069
rect 11060 23035 11112 23044
rect 11060 23001 11069 23035
rect 11069 23001 11103 23035
rect 11103 23001 11112 23035
rect 11060 22992 11112 23001
rect 11152 22992 11204 23044
rect 14004 22992 14056 23044
rect 14464 23035 14516 23044
rect 14464 23001 14473 23035
rect 14473 23001 14507 23035
rect 14507 23001 14516 23035
rect 14464 22992 14516 23001
rect 14648 22992 14700 23044
rect 7656 22924 7708 22976
rect 12532 22924 12584 22976
rect 13452 22924 13504 22976
rect 15844 23060 15896 23112
rect 17960 23128 18012 23180
rect 17132 23103 17184 23112
rect 17132 23069 17141 23103
rect 17141 23069 17175 23103
rect 17175 23069 17184 23103
rect 17132 23060 17184 23069
rect 17408 23103 17460 23112
rect 17408 23069 17417 23103
rect 17417 23069 17451 23103
rect 17451 23069 17460 23103
rect 17408 23060 17460 23069
rect 17684 23103 17736 23112
rect 17684 23069 17693 23103
rect 17693 23069 17727 23103
rect 17727 23069 17736 23103
rect 17684 23060 17736 23069
rect 17868 23060 17920 23112
rect 17316 22992 17368 23044
rect 17776 22992 17828 23044
rect 20536 23171 20588 23180
rect 20536 23137 20545 23171
rect 20545 23137 20579 23171
rect 20579 23137 20588 23171
rect 20536 23128 20588 23137
rect 22560 23264 22612 23316
rect 23296 23264 23348 23316
rect 23388 23264 23440 23316
rect 26056 23264 26108 23316
rect 26332 23264 26384 23316
rect 29368 23264 29420 23316
rect 32036 23264 32088 23316
rect 33048 23264 33100 23316
rect 34612 23264 34664 23316
rect 23480 23239 23532 23248
rect 23480 23205 23489 23239
rect 23489 23205 23523 23239
rect 23523 23205 23532 23239
rect 23480 23196 23532 23205
rect 27528 23196 27580 23248
rect 22192 23128 22244 23180
rect 23848 23128 23900 23180
rect 24860 23128 24912 23180
rect 18604 23103 18656 23112
rect 18604 23069 18613 23103
rect 18613 23069 18647 23103
rect 18647 23069 18656 23103
rect 20444 23103 20496 23112
rect 18604 23060 18656 23069
rect 20444 23069 20453 23103
rect 20453 23069 20487 23103
rect 20487 23069 20496 23103
rect 20444 23060 20496 23069
rect 20628 23060 20680 23112
rect 22284 23060 22336 23112
rect 22928 23103 22980 23112
rect 22928 23069 22937 23103
rect 22937 23069 22971 23103
rect 22971 23069 22980 23103
rect 22928 23060 22980 23069
rect 23020 23060 23072 23112
rect 15568 22924 15620 22976
rect 17500 22924 17552 22976
rect 19708 22992 19760 23044
rect 20260 22992 20312 23044
rect 22468 22992 22520 23044
rect 24032 23060 24084 23112
rect 24400 23060 24452 23112
rect 25136 23060 25188 23112
rect 24124 22992 24176 23044
rect 18788 22924 18840 22976
rect 23664 22924 23716 22976
rect 26056 23103 26108 23112
rect 26056 23069 26065 23103
rect 26065 23069 26099 23103
rect 26099 23069 26108 23103
rect 26056 23060 26108 23069
rect 27344 23060 27396 23112
rect 29736 23103 29788 23112
rect 29736 23069 29745 23103
rect 29745 23069 29779 23103
rect 29779 23069 29788 23103
rect 29736 23060 29788 23069
rect 29920 23103 29972 23112
rect 29920 23069 29929 23103
rect 29929 23069 29963 23103
rect 29963 23069 29972 23103
rect 29920 23060 29972 23069
rect 32404 23060 32456 23112
rect 32496 23103 32548 23112
rect 32496 23069 32505 23103
rect 32505 23069 32539 23103
rect 32539 23069 32548 23103
rect 32496 23060 32548 23069
rect 25872 23035 25924 23044
rect 25872 23001 25881 23035
rect 25881 23001 25915 23035
rect 25915 23001 25924 23035
rect 25872 22992 25924 23001
rect 25964 23035 26016 23044
rect 25964 23001 25973 23035
rect 25973 23001 26007 23035
rect 26007 23001 26016 23035
rect 25964 22992 26016 23001
rect 30012 23035 30064 23044
rect 30012 23001 30021 23035
rect 30021 23001 30055 23035
rect 30055 23001 30064 23035
rect 30012 22992 30064 23001
rect 32956 23060 33008 23112
rect 33324 22992 33376 23044
rect 34980 23103 35032 23112
rect 34980 23069 34989 23103
rect 34989 23069 35023 23103
rect 35023 23069 35032 23103
rect 34980 23060 35032 23069
rect 35072 23060 35124 23112
rect 35808 23128 35860 23180
rect 25688 22924 25740 22976
rect 26240 22967 26292 22976
rect 26240 22933 26249 22967
rect 26249 22933 26283 22967
rect 26283 22933 26292 22967
rect 26240 22924 26292 22933
rect 31852 22924 31904 22976
rect 32588 22924 32640 22976
rect 34336 22924 34388 22976
rect 36084 22967 36136 22976
rect 36084 22933 36093 22967
rect 36093 22933 36127 22967
rect 36127 22933 36136 22967
rect 36084 22924 36136 22933
rect 36176 22924 36228 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 2688 22720 2740 22772
rect 3148 22720 3200 22772
rect 3976 22763 4028 22772
rect 3976 22729 3985 22763
rect 3985 22729 4019 22763
rect 4019 22729 4028 22763
rect 3976 22720 4028 22729
rect 4436 22720 4488 22772
rect 2504 22652 2556 22704
rect 3056 22652 3108 22704
rect 4528 22652 4580 22704
rect 4804 22652 4856 22704
rect 5632 22720 5684 22772
rect 2964 22627 3016 22636
rect 2964 22593 2973 22627
rect 2973 22593 3007 22627
rect 3007 22593 3016 22627
rect 2964 22584 3016 22593
rect 3884 22627 3936 22636
rect 3884 22593 3893 22627
rect 3893 22593 3927 22627
rect 3927 22593 3936 22627
rect 3884 22584 3936 22593
rect 4068 22627 4120 22636
rect 4068 22593 4077 22627
rect 4077 22593 4111 22627
rect 4111 22593 4120 22627
rect 4068 22584 4120 22593
rect 4712 22584 4764 22636
rect 5172 22584 5224 22636
rect 2872 22516 2924 22568
rect 4896 22516 4948 22568
rect 5356 22516 5408 22568
rect 5908 22652 5960 22704
rect 7012 22720 7064 22772
rect 9128 22720 9180 22772
rect 9404 22720 9456 22772
rect 9864 22720 9916 22772
rect 11060 22763 11112 22772
rect 11060 22729 11069 22763
rect 11069 22729 11103 22763
rect 11103 22729 11112 22763
rect 11060 22720 11112 22729
rect 7380 22652 7432 22704
rect 7656 22652 7708 22704
rect 7932 22652 7984 22704
rect 11336 22652 11388 22704
rect 6920 22584 6972 22636
rect 8116 22584 8168 22636
rect 8760 22584 8812 22636
rect 3608 22448 3660 22500
rect 6276 22448 6328 22500
rect 10140 22584 10192 22636
rect 12348 22720 12400 22772
rect 12440 22720 12492 22772
rect 14096 22720 14148 22772
rect 15200 22720 15252 22772
rect 15476 22763 15528 22772
rect 15476 22729 15485 22763
rect 15485 22729 15519 22763
rect 15519 22729 15528 22763
rect 15476 22720 15528 22729
rect 15844 22720 15896 22772
rect 18512 22720 18564 22772
rect 20444 22763 20496 22772
rect 20444 22729 20453 22763
rect 20453 22729 20487 22763
rect 20487 22729 20496 22763
rect 20444 22720 20496 22729
rect 22928 22720 22980 22772
rect 14004 22652 14056 22704
rect 10048 22516 10100 22568
rect 11980 22559 12032 22568
rect 11980 22525 11989 22559
rect 11989 22525 12023 22559
rect 12023 22525 12032 22559
rect 11980 22516 12032 22525
rect 12164 22559 12216 22568
rect 12164 22525 12173 22559
rect 12173 22525 12207 22559
rect 12207 22525 12216 22559
rect 12164 22516 12216 22525
rect 3700 22380 3752 22432
rect 4160 22380 4212 22432
rect 6184 22380 6236 22432
rect 12440 22584 12492 22636
rect 12532 22627 12584 22636
rect 12532 22593 12541 22627
rect 12541 22593 12575 22627
rect 12575 22593 12584 22627
rect 12532 22584 12584 22593
rect 12808 22516 12860 22568
rect 13452 22584 13504 22636
rect 14188 22584 14240 22636
rect 16120 22695 16172 22704
rect 16120 22661 16129 22695
rect 16129 22661 16163 22695
rect 16163 22661 16172 22695
rect 16120 22652 16172 22661
rect 16764 22652 16816 22704
rect 17500 22652 17552 22704
rect 19340 22652 19392 22704
rect 23664 22720 23716 22772
rect 23756 22720 23808 22772
rect 25596 22720 25648 22772
rect 26240 22720 26292 22772
rect 27528 22763 27580 22772
rect 27528 22729 27537 22763
rect 27537 22729 27571 22763
rect 27571 22729 27580 22763
rect 27528 22720 27580 22729
rect 28356 22720 28408 22772
rect 29920 22720 29972 22772
rect 32496 22720 32548 22772
rect 33048 22720 33100 22772
rect 35072 22720 35124 22772
rect 14464 22584 14516 22636
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 15568 22584 15620 22636
rect 16856 22584 16908 22636
rect 17132 22627 17184 22636
rect 17132 22593 17141 22627
rect 17141 22593 17175 22627
rect 17175 22593 17184 22627
rect 17132 22584 17184 22593
rect 17316 22627 17368 22636
rect 17316 22593 17325 22627
rect 17325 22593 17359 22627
rect 17359 22593 17368 22627
rect 17316 22584 17368 22593
rect 17868 22627 17920 22636
rect 17868 22593 17877 22627
rect 17877 22593 17911 22627
rect 17911 22593 17920 22627
rect 17868 22584 17920 22593
rect 20720 22627 20772 22636
rect 20720 22593 20729 22627
rect 20729 22593 20763 22627
rect 20763 22593 20772 22627
rect 20720 22584 20772 22593
rect 21916 22584 21968 22636
rect 22192 22627 22244 22636
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 22468 22584 22520 22636
rect 14188 22380 14240 22432
rect 16304 22516 16356 22568
rect 17500 22516 17552 22568
rect 23296 22584 23348 22636
rect 23388 22627 23440 22636
rect 23388 22593 23397 22627
rect 23397 22593 23431 22627
rect 23431 22593 23440 22627
rect 23388 22584 23440 22593
rect 23572 22627 23624 22636
rect 23572 22593 23581 22627
rect 23581 22593 23615 22627
rect 23615 22593 23624 22627
rect 23572 22584 23624 22593
rect 24032 22627 24084 22636
rect 24032 22593 24041 22627
rect 24041 22593 24075 22627
rect 24075 22593 24084 22627
rect 24032 22584 24084 22593
rect 16028 22448 16080 22500
rect 16764 22448 16816 22500
rect 19248 22448 19300 22500
rect 20076 22448 20128 22500
rect 21824 22380 21876 22432
rect 24124 22516 24176 22568
rect 25780 22627 25832 22636
rect 25780 22593 25789 22627
rect 25789 22593 25823 22627
rect 25823 22593 25832 22627
rect 25780 22584 25832 22593
rect 26148 22584 26200 22636
rect 26516 22584 26568 22636
rect 26608 22584 26660 22636
rect 27160 22627 27212 22636
rect 27160 22593 27169 22627
rect 27169 22593 27203 22627
rect 27203 22593 27212 22627
rect 27160 22584 27212 22593
rect 25872 22516 25924 22568
rect 23940 22491 23992 22500
rect 23940 22457 23949 22491
rect 23949 22457 23983 22491
rect 23983 22457 23992 22491
rect 23940 22448 23992 22457
rect 26056 22448 26108 22500
rect 27436 22584 27488 22636
rect 27712 22627 27764 22636
rect 27712 22593 27721 22627
rect 27721 22593 27755 22627
rect 27755 22593 27764 22627
rect 27712 22584 27764 22593
rect 30196 22627 30248 22636
rect 30196 22593 30205 22627
rect 30205 22593 30239 22627
rect 30239 22593 30248 22627
rect 30196 22584 30248 22593
rect 32128 22627 32180 22636
rect 32128 22593 32137 22627
rect 32137 22593 32171 22627
rect 32171 22593 32180 22627
rect 32128 22584 32180 22593
rect 32404 22584 32456 22636
rect 33048 22584 33100 22636
rect 36176 22652 36228 22704
rect 36452 22720 36504 22772
rect 33232 22627 33284 22636
rect 33232 22593 33241 22627
rect 33241 22593 33275 22627
rect 33275 22593 33284 22627
rect 33232 22584 33284 22593
rect 33324 22584 33376 22636
rect 34428 22584 34480 22636
rect 34980 22584 35032 22636
rect 35348 22627 35400 22636
rect 35348 22593 35357 22627
rect 35357 22593 35391 22627
rect 35391 22593 35400 22627
rect 35348 22584 35400 22593
rect 35808 22584 35860 22636
rect 31852 22516 31904 22568
rect 32956 22559 33008 22568
rect 32956 22525 32965 22559
rect 32965 22525 32999 22559
rect 32999 22525 33008 22559
rect 32956 22516 33008 22525
rect 36268 22627 36320 22636
rect 36268 22593 36277 22627
rect 36277 22593 36311 22627
rect 36311 22593 36320 22627
rect 36268 22584 36320 22593
rect 33232 22448 33284 22500
rect 37556 22584 37608 22636
rect 37832 22491 37884 22500
rect 37832 22457 37841 22491
rect 37841 22457 37875 22491
rect 37875 22457 37884 22491
rect 37832 22448 37884 22457
rect 24768 22380 24820 22432
rect 25964 22380 26016 22432
rect 29736 22380 29788 22432
rect 30656 22423 30708 22432
rect 30656 22389 30665 22423
rect 30665 22389 30699 22423
rect 30699 22389 30708 22423
rect 30656 22380 30708 22389
rect 32496 22423 32548 22432
rect 32496 22389 32505 22423
rect 32505 22389 32539 22423
rect 32539 22389 32548 22423
rect 32496 22380 32548 22389
rect 32588 22380 32640 22432
rect 34796 22380 34848 22432
rect 35900 22380 35952 22432
rect 36452 22423 36504 22432
rect 36452 22389 36461 22423
rect 36461 22389 36495 22423
rect 36495 22389 36504 22423
rect 36452 22380 36504 22389
rect 37004 22423 37056 22432
rect 37004 22389 37013 22423
rect 37013 22389 37047 22423
rect 37047 22389 37056 22423
rect 37004 22380 37056 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3608 22176 3660 22228
rect 9680 22176 9732 22228
rect 11980 22176 12032 22228
rect 1952 22015 2004 22024
rect 1952 21981 1961 22015
rect 1961 21981 1995 22015
rect 1995 21981 2004 22015
rect 1952 21972 2004 21981
rect 4068 21972 4120 22024
rect 6000 22108 6052 22160
rect 6276 22108 6328 22160
rect 25872 22176 25924 22228
rect 15384 22108 15436 22160
rect 16396 22108 16448 22160
rect 16764 22108 16816 22160
rect 10048 22083 10100 22092
rect 10048 22049 10057 22083
rect 10057 22049 10091 22083
rect 10091 22049 10100 22083
rect 10048 22040 10100 22049
rect 3884 21904 3936 21956
rect 11428 21972 11480 22024
rect 12164 22040 12216 22092
rect 14372 22040 14424 22092
rect 15660 22040 15712 22092
rect 13728 21972 13780 22024
rect 14188 21972 14240 22024
rect 1768 21879 1820 21888
rect 1768 21845 1777 21879
rect 1777 21845 1811 21879
rect 1811 21845 1820 21879
rect 1768 21836 1820 21845
rect 14556 21904 14608 21956
rect 15384 21972 15436 22024
rect 15476 22015 15528 22024
rect 15476 21981 15485 22015
rect 15485 21981 15519 22015
rect 15519 21981 15528 22015
rect 15476 21972 15528 21981
rect 15568 22015 15620 22024
rect 15568 21981 15577 22015
rect 15577 21981 15611 22015
rect 15611 21981 15620 22015
rect 15568 21972 15620 21981
rect 16948 22108 17000 22160
rect 17224 22108 17276 22160
rect 17868 22108 17920 22160
rect 19248 22151 19300 22160
rect 19248 22117 19257 22151
rect 19257 22117 19291 22151
rect 19291 22117 19300 22151
rect 19248 22108 19300 22117
rect 23572 22108 23624 22160
rect 24584 22108 24636 22160
rect 24952 22108 25004 22160
rect 16120 21972 16172 22024
rect 16304 21972 16356 22024
rect 16396 22015 16448 22024
rect 16396 21981 16405 22015
rect 16405 21981 16439 22015
rect 16439 21981 16448 22015
rect 16396 21972 16448 21981
rect 16764 21972 16816 22024
rect 15108 21904 15160 21956
rect 17040 22015 17092 22024
rect 17040 21981 17049 22015
rect 17049 21981 17083 22015
rect 17083 21981 17092 22015
rect 17040 21972 17092 21981
rect 17132 21972 17184 22024
rect 19248 21972 19300 22024
rect 16948 21904 17000 21956
rect 19340 21904 19392 21956
rect 4344 21879 4396 21888
rect 4344 21845 4353 21879
rect 4353 21845 4387 21879
rect 4387 21845 4396 21879
rect 4344 21836 4396 21845
rect 5816 21836 5868 21888
rect 6920 21836 6972 21888
rect 8116 21836 8168 21888
rect 8484 21836 8536 21888
rect 9772 21879 9824 21888
rect 9772 21845 9781 21879
rect 9781 21845 9815 21879
rect 9815 21845 9824 21879
rect 9772 21836 9824 21845
rect 10876 21836 10928 21888
rect 11704 21879 11756 21888
rect 11704 21845 11713 21879
rect 11713 21845 11747 21879
rect 11747 21845 11756 21879
rect 11704 21836 11756 21845
rect 11796 21879 11848 21888
rect 11796 21845 11805 21879
rect 11805 21845 11839 21879
rect 11839 21845 11848 21879
rect 11796 21836 11848 21845
rect 12164 21836 12216 21888
rect 12992 21836 13044 21888
rect 16212 21836 16264 21888
rect 17592 21836 17644 21888
rect 19432 21836 19484 21888
rect 19984 22015 20036 22024
rect 19984 21981 19993 22015
rect 19993 21981 20027 22015
rect 20027 21981 20036 22015
rect 19984 21972 20036 21981
rect 20168 22015 20220 22024
rect 20168 21981 20177 22015
rect 20177 21981 20211 22015
rect 20211 21981 20220 22015
rect 20168 21972 20220 21981
rect 22008 21972 22060 22024
rect 22284 21972 22336 22024
rect 23480 21972 23532 22024
rect 24032 22040 24084 22092
rect 24492 21972 24544 22024
rect 24768 21972 24820 22024
rect 25320 22083 25372 22092
rect 25320 22049 25329 22083
rect 25329 22049 25363 22083
rect 25363 22049 25372 22083
rect 25320 22040 25372 22049
rect 26056 22040 26108 22092
rect 26608 22040 26660 22092
rect 19892 21904 19944 21956
rect 20352 21904 20404 21956
rect 23020 21904 23072 21956
rect 23388 21904 23440 21956
rect 25688 21972 25740 22024
rect 25780 22015 25832 22024
rect 25780 21981 25789 22015
rect 25789 21981 25823 22015
rect 25823 21981 25832 22015
rect 25780 21972 25832 21981
rect 26240 22015 26292 22024
rect 26240 21981 26243 22015
rect 26243 21981 26292 22015
rect 26240 21972 26292 21981
rect 26516 21972 26568 22024
rect 28264 22176 28316 22228
rect 28448 22176 28500 22228
rect 27528 22040 27580 22092
rect 22100 21836 22152 21888
rect 22468 21836 22520 21888
rect 28448 21972 28500 22024
rect 28724 21972 28776 22024
rect 30012 22040 30064 22092
rect 29092 21972 29144 22024
rect 31024 22108 31076 22160
rect 30564 21972 30616 22024
rect 31944 22108 31996 22160
rect 31852 22015 31904 22024
rect 31852 21981 31861 22015
rect 31861 21981 31895 22015
rect 31895 21981 31904 22015
rect 31852 21972 31904 21981
rect 32036 21972 32088 22024
rect 32772 22108 32824 22160
rect 33232 22176 33284 22228
rect 33324 22176 33376 22228
rect 33232 22083 33284 22092
rect 33232 22049 33241 22083
rect 33241 22049 33275 22083
rect 33275 22049 33284 22083
rect 33232 22040 33284 22049
rect 33508 22040 33560 22092
rect 35624 22040 35676 22092
rect 36176 22176 36228 22228
rect 36084 22040 36136 22092
rect 27528 21836 27580 21888
rect 27620 21879 27672 21888
rect 27620 21845 27629 21879
rect 27629 21845 27663 21879
rect 27663 21845 27672 21879
rect 27620 21836 27672 21845
rect 27712 21836 27764 21888
rect 27804 21836 27856 21888
rect 28264 21947 28316 21956
rect 28264 21913 28273 21947
rect 28273 21913 28307 21947
rect 28307 21913 28316 21947
rect 28264 21904 28316 21913
rect 28540 21879 28592 21888
rect 28540 21845 28549 21879
rect 28549 21845 28583 21879
rect 28583 21845 28592 21879
rect 28540 21836 28592 21845
rect 29000 21836 29052 21888
rect 31116 21947 31168 21956
rect 31116 21913 31125 21947
rect 31125 21913 31159 21947
rect 31159 21913 31168 21947
rect 31116 21904 31168 21913
rect 30380 21836 30432 21888
rect 30472 21836 30524 21888
rect 32680 22015 32732 22024
rect 32680 21981 32689 22015
rect 32689 21981 32723 22015
rect 32723 21981 32732 22015
rect 32680 21972 32732 21981
rect 34428 21972 34480 22024
rect 34796 21972 34848 22024
rect 35256 21972 35308 22024
rect 32588 21904 32640 21956
rect 34704 21879 34756 21888
rect 34704 21845 34713 21879
rect 34713 21845 34747 21879
rect 34747 21845 34756 21879
rect 34704 21836 34756 21845
rect 35716 21836 35768 21888
rect 36452 22040 36504 22092
rect 36912 21972 36964 22024
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 1768 21632 1820 21684
rect 1952 21632 2004 21684
rect 4344 21632 4396 21684
rect 2780 21496 2832 21548
rect 3608 21539 3660 21548
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 4712 21632 4764 21684
rect 5172 21607 5224 21616
rect 5172 21573 5181 21607
rect 5181 21573 5215 21607
rect 5215 21573 5224 21607
rect 5172 21564 5224 21573
rect 6920 21564 6972 21616
rect 7288 21564 7340 21616
rect 3056 21292 3108 21344
rect 5724 21539 5776 21548
rect 5724 21505 5733 21539
rect 5733 21505 5767 21539
rect 5767 21505 5776 21539
rect 5724 21496 5776 21505
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 5816 21496 5868 21505
rect 6184 21496 6236 21548
rect 4620 21360 4672 21412
rect 5080 21360 5132 21412
rect 6828 21471 6880 21480
rect 6828 21437 6837 21471
rect 6837 21437 6871 21471
rect 6871 21437 6880 21471
rect 6828 21428 6880 21437
rect 8852 21632 8904 21684
rect 9312 21632 9364 21684
rect 11244 21632 11296 21684
rect 14740 21632 14792 21684
rect 14924 21675 14976 21684
rect 14924 21641 14933 21675
rect 14933 21641 14967 21675
rect 14967 21641 14976 21675
rect 14924 21632 14976 21641
rect 8576 21496 8628 21548
rect 9680 21539 9732 21548
rect 9680 21505 9689 21539
rect 9689 21505 9723 21539
rect 9723 21505 9732 21539
rect 9680 21496 9732 21505
rect 9864 21496 9916 21548
rect 9956 21539 10008 21548
rect 9956 21505 9965 21539
rect 9965 21505 9999 21539
rect 9999 21505 10008 21539
rect 9956 21496 10008 21505
rect 10048 21539 10100 21548
rect 10048 21505 10057 21539
rect 10057 21505 10091 21539
rect 10091 21505 10100 21539
rect 10048 21496 10100 21505
rect 10324 21539 10376 21548
rect 10324 21505 10333 21539
rect 10333 21505 10367 21539
rect 10367 21505 10376 21539
rect 10324 21496 10376 21505
rect 12440 21496 12492 21548
rect 13360 21496 13412 21548
rect 13912 21564 13964 21616
rect 14004 21564 14056 21616
rect 14096 21496 14148 21548
rect 14188 21496 14240 21548
rect 11980 21471 12032 21480
rect 11980 21437 11989 21471
rect 11989 21437 12023 21471
rect 12023 21437 12032 21471
rect 11980 21428 12032 21437
rect 12164 21471 12216 21480
rect 12164 21437 12173 21471
rect 12173 21437 12207 21471
rect 12207 21437 12216 21471
rect 12164 21428 12216 21437
rect 13636 21471 13688 21480
rect 13636 21437 13645 21471
rect 13645 21437 13679 21471
rect 13679 21437 13688 21471
rect 13636 21428 13688 21437
rect 14372 21496 14424 21548
rect 17132 21632 17184 21684
rect 17408 21632 17460 21684
rect 17500 21632 17552 21684
rect 18972 21675 19024 21684
rect 18972 21641 18981 21675
rect 18981 21641 19015 21675
rect 19015 21641 19024 21675
rect 18972 21632 19024 21641
rect 15200 21539 15252 21548
rect 15200 21505 15209 21539
rect 15209 21505 15243 21539
rect 15243 21505 15252 21539
rect 15200 21496 15252 21505
rect 15292 21539 15344 21548
rect 15292 21505 15301 21539
rect 15301 21505 15335 21539
rect 15335 21505 15344 21539
rect 15292 21496 15344 21505
rect 15384 21496 15436 21548
rect 15936 21564 15988 21616
rect 16304 21564 16356 21616
rect 16580 21564 16632 21616
rect 20076 21632 20128 21684
rect 20168 21675 20220 21684
rect 20168 21641 20177 21675
rect 20177 21641 20211 21675
rect 20211 21641 20220 21675
rect 20168 21632 20220 21641
rect 20352 21632 20404 21684
rect 22192 21632 22244 21684
rect 24676 21632 24728 21684
rect 19340 21564 19392 21616
rect 16948 21496 17000 21548
rect 17132 21496 17184 21548
rect 17960 21496 18012 21548
rect 19248 21496 19300 21548
rect 18052 21471 18104 21480
rect 18052 21437 18061 21471
rect 18061 21437 18095 21471
rect 18095 21437 18104 21471
rect 18052 21428 18104 21437
rect 18144 21471 18196 21480
rect 18144 21437 18153 21471
rect 18153 21437 18187 21471
rect 18187 21437 18196 21471
rect 18144 21428 18196 21437
rect 18972 21428 19024 21480
rect 19432 21471 19484 21480
rect 19432 21437 19441 21471
rect 19441 21437 19475 21471
rect 19475 21437 19484 21471
rect 19432 21428 19484 21437
rect 21180 21564 21232 21616
rect 22008 21564 22060 21616
rect 23848 21564 23900 21616
rect 24768 21564 24820 21616
rect 25136 21632 25188 21684
rect 26700 21632 26752 21684
rect 27712 21675 27764 21684
rect 27712 21641 27721 21675
rect 27721 21641 27755 21675
rect 27755 21641 27764 21675
rect 27712 21632 27764 21641
rect 29920 21675 29972 21684
rect 29920 21641 29929 21675
rect 29929 21641 29963 21675
rect 29963 21641 29972 21675
rect 29920 21632 29972 21641
rect 30380 21632 30432 21684
rect 32588 21675 32640 21684
rect 32588 21641 32597 21675
rect 32597 21641 32631 21675
rect 32631 21641 32640 21675
rect 32588 21632 32640 21641
rect 25320 21564 25372 21616
rect 25872 21564 25924 21616
rect 20352 21539 20404 21548
rect 20352 21505 20361 21539
rect 20361 21505 20395 21539
rect 20395 21505 20404 21539
rect 20352 21496 20404 21505
rect 19984 21428 20036 21480
rect 8300 21403 8352 21412
rect 8300 21369 8309 21403
rect 8309 21369 8343 21403
rect 8343 21369 8352 21403
rect 8300 21360 8352 21369
rect 16580 21360 16632 21412
rect 4896 21292 4948 21344
rect 6644 21292 6696 21344
rect 8116 21292 8168 21344
rect 10968 21292 11020 21344
rect 22928 21360 22980 21412
rect 23296 21428 23348 21480
rect 17132 21292 17184 21344
rect 23480 21360 23532 21412
rect 25136 21539 25188 21548
rect 25136 21505 25145 21539
rect 25145 21505 25179 21539
rect 25179 21505 25188 21539
rect 25136 21496 25188 21505
rect 25504 21496 25556 21548
rect 26056 21496 26108 21548
rect 27896 21564 27948 21616
rect 28816 21564 28868 21616
rect 29736 21607 29788 21616
rect 29736 21573 29745 21607
rect 29745 21573 29779 21607
rect 29779 21573 29788 21607
rect 29736 21564 29788 21573
rect 27712 21539 27764 21548
rect 27712 21505 27721 21539
rect 27721 21505 27755 21539
rect 27755 21505 27764 21539
rect 27712 21496 27764 21505
rect 30564 21496 30616 21548
rect 33784 21632 33836 21684
rect 34704 21632 34756 21684
rect 35256 21675 35308 21684
rect 35256 21641 35265 21675
rect 35265 21641 35299 21675
rect 35299 21641 35308 21675
rect 35256 21632 35308 21641
rect 31116 21496 31168 21548
rect 31944 21496 31996 21548
rect 32680 21539 32732 21548
rect 32680 21505 32689 21539
rect 32689 21505 32723 21539
rect 32723 21505 32732 21539
rect 32680 21496 32732 21505
rect 33324 21539 33376 21548
rect 33324 21505 33333 21539
rect 33333 21505 33367 21539
rect 33367 21505 33376 21539
rect 33324 21496 33376 21505
rect 33600 21496 33652 21548
rect 33784 21539 33836 21548
rect 33784 21505 33793 21539
rect 33793 21505 33827 21539
rect 33827 21505 33836 21539
rect 33784 21496 33836 21505
rect 35348 21564 35400 21616
rect 35716 21496 35768 21548
rect 35808 21539 35860 21548
rect 35808 21505 35817 21539
rect 35817 21505 35851 21539
rect 35851 21505 35860 21539
rect 35808 21496 35860 21505
rect 36176 21496 36228 21548
rect 36452 21496 36504 21548
rect 27436 21360 27488 21412
rect 28724 21360 28776 21412
rect 35624 21428 35676 21480
rect 37188 21428 37240 21480
rect 23112 21335 23164 21344
rect 23112 21301 23121 21335
rect 23121 21301 23155 21335
rect 23155 21301 23164 21335
rect 23112 21292 23164 21301
rect 29184 21292 29236 21344
rect 29644 21292 29696 21344
rect 30932 21335 30984 21344
rect 30932 21301 30941 21335
rect 30941 21301 30975 21335
rect 30975 21301 30984 21335
rect 30932 21292 30984 21301
rect 33232 21292 33284 21344
rect 35440 21335 35492 21344
rect 35440 21301 35449 21335
rect 35449 21301 35483 21335
rect 35483 21301 35492 21335
rect 35440 21292 35492 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 4620 21088 4672 21140
rect 6828 21088 6880 21140
rect 4068 20995 4120 21004
rect 4068 20961 4077 20995
rect 4077 20961 4111 20995
rect 4111 20961 4120 20995
rect 4068 20952 4120 20961
rect 1860 20884 1912 20936
rect 3516 20884 3568 20936
rect 3608 20884 3660 20936
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 6920 20884 6972 20936
rect 8300 21088 8352 21140
rect 9772 21088 9824 21140
rect 10140 21131 10192 21140
rect 10140 21097 10149 21131
rect 10149 21097 10183 21131
rect 10183 21097 10192 21131
rect 10140 21088 10192 21097
rect 12164 21088 12216 21140
rect 7932 20952 7984 21004
rect 14004 21020 14056 21072
rect 14740 21088 14792 21140
rect 15476 21131 15528 21140
rect 15476 21097 15485 21131
rect 15485 21097 15519 21131
rect 15519 21097 15528 21131
rect 15476 21088 15528 21097
rect 17040 21088 17092 21140
rect 17132 21088 17184 21140
rect 18236 21088 18288 21140
rect 18512 21088 18564 21140
rect 18788 21088 18840 21140
rect 17500 21020 17552 21072
rect 20352 21088 20404 21140
rect 21088 21088 21140 21140
rect 21824 21088 21876 21140
rect 25044 21131 25096 21140
rect 25044 21097 25053 21131
rect 25053 21097 25087 21131
rect 25087 21097 25096 21131
rect 25044 21088 25096 21097
rect 25320 21088 25372 21140
rect 26976 21088 27028 21140
rect 27528 21088 27580 21140
rect 30932 21088 30984 21140
rect 33508 21088 33560 21140
rect 35256 21088 35308 21140
rect 35440 21088 35492 21140
rect 8668 20884 8720 20936
rect 10048 20952 10100 21004
rect 12348 20952 12400 21004
rect 9588 20927 9640 20936
rect 9588 20893 9597 20927
rect 9597 20893 9631 20927
rect 9631 20893 9640 20927
rect 9588 20884 9640 20893
rect 9956 20927 10008 20936
rect 9956 20893 9965 20927
rect 9965 20893 9999 20927
rect 9999 20893 10008 20927
rect 9956 20884 10008 20893
rect 13912 20884 13964 20936
rect 14188 20884 14240 20936
rect 20904 20952 20956 21004
rect 21916 21020 21968 21072
rect 23112 21020 23164 21072
rect 1492 20791 1544 20800
rect 1492 20757 1501 20791
rect 1501 20757 1535 20791
rect 1535 20757 1544 20791
rect 1492 20748 1544 20757
rect 2872 20748 2924 20800
rect 4068 20748 4120 20800
rect 5632 20859 5684 20868
rect 5632 20825 5641 20859
rect 5641 20825 5675 20859
rect 5675 20825 5684 20859
rect 5632 20816 5684 20825
rect 9220 20859 9272 20868
rect 9220 20825 9229 20859
rect 9229 20825 9263 20859
rect 9263 20825 9272 20859
rect 9220 20816 9272 20825
rect 9772 20859 9824 20868
rect 9772 20825 9781 20859
rect 9781 20825 9815 20859
rect 9815 20825 9824 20859
rect 9772 20816 9824 20825
rect 9864 20859 9916 20868
rect 9864 20825 9873 20859
rect 9873 20825 9907 20859
rect 9907 20825 9916 20859
rect 9864 20816 9916 20825
rect 10600 20816 10652 20868
rect 14004 20816 14056 20868
rect 11428 20748 11480 20800
rect 12808 20748 12860 20800
rect 14096 20748 14148 20800
rect 14924 20859 14976 20868
rect 14924 20825 14933 20859
rect 14933 20825 14967 20859
rect 14967 20825 14976 20859
rect 14924 20816 14976 20825
rect 17132 20927 17184 20936
rect 17132 20893 17136 20927
rect 17136 20893 17170 20927
rect 17170 20893 17184 20927
rect 17132 20884 17184 20893
rect 17868 20884 17920 20936
rect 18788 20884 18840 20936
rect 14556 20748 14608 20800
rect 15200 20748 15252 20800
rect 15476 20748 15528 20800
rect 15660 20748 15712 20800
rect 17408 20816 17460 20868
rect 17592 20748 17644 20800
rect 18512 20748 18564 20800
rect 19984 20884 20036 20936
rect 20352 20927 20404 20936
rect 20352 20893 20361 20927
rect 20361 20893 20395 20927
rect 20395 20893 20404 20927
rect 20352 20884 20404 20893
rect 20444 20884 20496 20936
rect 20812 20927 20864 20936
rect 20812 20893 20821 20927
rect 20821 20893 20855 20927
rect 20855 20893 20864 20927
rect 20812 20884 20864 20893
rect 22100 20952 22152 21004
rect 21180 20884 21232 20936
rect 21456 20927 21508 20936
rect 21456 20893 21466 20927
rect 21466 20893 21500 20927
rect 21500 20893 21508 20927
rect 21456 20884 21508 20893
rect 21824 20927 21876 20936
rect 21824 20893 21838 20927
rect 21838 20893 21872 20927
rect 21872 20893 21876 20927
rect 21824 20884 21876 20893
rect 22192 20927 22244 20936
rect 22192 20893 22201 20927
rect 22201 20893 22235 20927
rect 22235 20893 22244 20927
rect 22192 20884 22244 20893
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 22928 20952 22980 21004
rect 23388 20952 23440 21004
rect 24952 20952 25004 21004
rect 24400 20884 24452 20936
rect 24860 20884 24912 20936
rect 25504 21020 25556 21072
rect 25688 21020 25740 21072
rect 34336 21020 34388 21072
rect 19340 20748 19392 20800
rect 20352 20748 20404 20800
rect 20444 20748 20496 20800
rect 21088 20748 21140 20800
rect 22008 20791 22060 20800
rect 22008 20757 22017 20791
rect 22017 20757 22051 20791
rect 22051 20757 22060 20791
rect 22008 20748 22060 20757
rect 22192 20748 22244 20800
rect 24492 20816 24544 20868
rect 22836 20791 22888 20800
rect 22836 20757 22845 20791
rect 22845 20757 22879 20791
rect 22879 20757 22888 20791
rect 22836 20748 22888 20757
rect 24860 20791 24912 20800
rect 24860 20757 24869 20791
rect 24869 20757 24903 20791
rect 24903 20757 24912 20791
rect 24860 20748 24912 20757
rect 26700 20884 26752 20936
rect 27436 20952 27488 21004
rect 27252 20884 27304 20936
rect 30656 20995 30708 21004
rect 30656 20961 30665 20995
rect 30665 20961 30699 20995
rect 30699 20961 30708 20995
rect 30656 20952 30708 20961
rect 32312 20952 32364 21004
rect 33048 20952 33100 21004
rect 35348 21020 35400 21072
rect 29460 20884 29512 20936
rect 30380 20927 30432 20936
rect 30380 20893 30389 20927
rect 30389 20893 30423 20927
rect 30423 20893 30432 20927
rect 30380 20884 30432 20893
rect 30472 20884 30524 20936
rect 33416 20884 33468 20936
rect 26884 20816 26936 20868
rect 27620 20748 27672 20800
rect 30196 20791 30248 20800
rect 30196 20757 30205 20791
rect 30205 20757 30239 20791
rect 30239 20757 30248 20791
rect 30196 20748 30248 20757
rect 33324 20816 33376 20868
rect 35256 20884 35308 20936
rect 35440 20927 35492 20936
rect 35440 20893 35449 20927
rect 35449 20893 35483 20927
rect 35483 20893 35492 20927
rect 35440 20884 35492 20893
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 38384 20680 38436 20732
rect 3148 20408 3200 20460
rect 2872 20383 2924 20392
rect 2872 20349 2881 20383
rect 2881 20349 2915 20383
rect 2915 20349 2924 20383
rect 2872 20340 2924 20349
rect 3056 20383 3108 20392
rect 3056 20349 3065 20383
rect 3065 20349 3099 20383
rect 3099 20349 3108 20383
rect 3056 20340 3108 20349
rect 3608 20408 3660 20460
rect 3884 20544 3936 20596
rect 13176 20544 13228 20596
rect 14280 20544 14332 20596
rect 15568 20544 15620 20596
rect 15660 20587 15712 20596
rect 15660 20553 15669 20587
rect 15669 20553 15703 20587
rect 15703 20553 15712 20587
rect 15660 20544 15712 20553
rect 9772 20476 9824 20528
rect 14004 20476 14056 20528
rect 3976 20408 4028 20460
rect 11980 20408 12032 20460
rect 14648 20519 14700 20528
rect 14648 20485 14657 20519
rect 14657 20485 14691 20519
rect 14691 20485 14700 20519
rect 14648 20476 14700 20485
rect 15108 20476 15160 20528
rect 16120 20544 16172 20596
rect 18604 20544 18656 20596
rect 18880 20544 18932 20596
rect 20444 20544 20496 20596
rect 21088 20544 21140 20596
rect 7380 20340 7432 20392
rect 7932 20340 7984 20392
rect 8392 20340 8444 20392
rect 11612 20383 11664 20392
rect 11612 20349 11621 20383
rect 11621 20349 11655 20383
rect 11655 20349 11664 20383
rect 11612 20340 11664 20349
rect 3792 20272 3844 20324
rect 12256 20272 12308 20324
rect 15568 20451 15620 20460
rect 15568 20417 15577 20451
rect 15577 20417 15611 20451
rect 15611 20417 15620 20451
rect 15568 20408 15620 20417
rect 15108 20340 15160 20392
rect 17776 20408 17828 20460
rect 17960 20408 18012 20460
rect 18144 20451 18196 20460
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 18144 20408 18196 20417
rect 18420 20408 18472 20460
rect 18512 20451 18564 20460
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 18604 20451 18656 20460
rect 18604 20417 18613 20451
rect 18613 20417 18647 20451
rect 18647 20417 18656 20451
rect 18604 20408 18656 20417
rect 19248 20451 19300 20460
rect 16120 20340 16172 20392
rect 16948 20340 17000 20392
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 20076 20451 20128 20460
rect 20076 20417 20085 20451
rect 20085 20417 20119 20451
rect 20119 20417 20128 20451
rect 20076 20408 20128 20417
rect 20352 20451 20404 20460
rect 20352 20417 20361 20451
rect 20361 20417 20395 20451
rect 20395 20417 20404 20451
rect 20352 20408 20404 20417
rect 19064 20340 19116 20392
rect 20628 20451 20680 20460
rect 20628 20417 20637 20451
rect 20637 20417 20671 20451
rect 20671 20417 20680 20451
rect 20628 20408 20680 20417
rect 20904 20451 20956 20460
rect 20904 20417 20913 20451
rect 20913 20417 20947 20451
rect 20947 20417 20956 20451
rect 20904 20408 20956 20417
rect 23296 20544 23348 20596
rect 23388 20544 23440 20596
rect 25504 20544 25556 20596
rect 27988 20544 28040 20596
rect 35808 20544 35860 20596
rect 32036 20476 32088 20528
rect 33324 20476 33376 20528
rect 22100 20340 22152 20392
rect 23572 20340 23624 20392
rect 18052 20272 18104 20324
rect 22284 20272 22336 20324
rect 24400 20451 24452 20460
rect 24400 20417 24409 20451
rect 24409 20417 24443 20451
rect 24443 20417 24452 20451
rect 24400 20408 24452 20417
rect 24584 20451 24636 20460
rect 24584 20417 24593 20451
rect 24593 20417 24627 20451
rect 24627 20417 24636 20451
rect 24584 20408 24636 20417
rect 24860 20408 24912 20460
rect 24676 20272 24728 20324
rect 25228 20408 25280 20460
rect 25872 20408 25924 20460
rect 26056 20451 26108 20460
rect 26056 20417 26065 20451
rect 26065 20417 26099 20451
rect 26099 20417 26108 20451
rect 26056 20408 26108 20417
rect 26240 20408 26292 20460
rect 26700 20408 26752 20460
rect 27252 20451 27304 20460
rect 27252 20417 27261 20451
rect 27261 20417 27295 20451
rect 27295 20417 27304 20451
rect 27252 20408 27304 20417
rect 25320 20383 25372 20392
rect 25320 20349 25329 20383
rect 25329 20349 25363 20383
rect 25363 20349 25372 20383
rect 25320 20340 25372 20349
rect 25412 20340 25464 20392
rect 26148 20272 26200 20324
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 3976 20204 4028 20256
rect 7196 20247 7248 20256
rect 7196 20213 7205 20247
rect 7205 20213 7239 20247
rect 7239 20213 7248 20247
rect 7196 20204 7248 20213
rect 11888 20204 11940 20256
rect 16304 20204 16356 20256
rect 17776 20204 17828 20256
rect 18604 20204 18656 20256
rect 19340 20204 19392 20256
rect 19892 20204 19944 20256
rect 20168 20204 20220 20256
rect 20352 20204 20404 20256
rect 21456 20204 21508 20256
rect 21916 20204 21968 20256
rect 24032 20204 24084 20256
rect 24124 20247 24176 20256
rect 24124 20213 24133 20247
rect 24133 20213 24167 20247
rect 24167 20213 24176 20247
rect 24124 20204 24176 20213
rect 24952 20247 25004 20256
rect 24952 20213 24961 20247
rect 24961 20213 24995 20247
rect 24995 20213 25004 20247
rect 24952 20204 25004 20213
rect 25504 20204 25556 20256
rect 27620 20451 27672 20460
rect 27620 20417 27629 20451
rect 27629 20417 27663 20451
rect 27663 20417 27672 20451
rect 27620 20408 27672 20417
rect 28724 20340 28776 20392
rect 28816 20340 28868 20392
rect 29552 20408 29604 20460
rect 30380 20408 30432 20460
rect 30656 20408 30708 20460
rect 30932 20408 30984 20460
rect 31116 20408 31168 20460
rect 32588 20408 32640 20460
rect 35900 20451 35952 20460
rect 35900 20417 35909 20451
rect 35909 20417 35943 20451
rect 35943 20417 35952 20451
rect 35900 20408 35952 20417
rect 29644 20383 29696 20392
rect 29644 20349 29653 20383
rect 29653 20349 29687 20383
rect 29687 20349 29696 20383
rect 29644 20340 29696 20349
rect 27252 20272 27304 20324
rect 27528 20272 27580 20324
rect 28632 20272 28684 20324
rect 30656 20315 30708 20324
rect 30656 20281 30665 20315
rect 30665 20281 30699 20315
rect 30699 20281 30708 20315
rect 30656 20272 30708 20281
rect 33232 20383 33284 20392
rect 33232 20349 33241 20383
rect 33241 20349 33275 20383
rect 33275 20349 33284 20383
rect 33232 20340 33284 20349
rect 34428 20340 34480 20392
rect 33140 20272 33192 20324
rect 34520 20272 34572 20324
rect 35808 20383 35860 20392
rect 35808 20349 35817 20383
rect 35817 20349 35851 20383
rect 35851 20349 35860 20383
rect 35808 20340 35860 20349
rect 28908 20247 28960 20256
rect 28908 20213 28917 20247
rect 28917 20213 28951 20247
rect 28951 20213 28960 20247
rect 28908 20204 28960 20213
rect 31208 20204 31260 20256
rect 34796 20204 34848 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2412 20000 2464 20052
rect 2872 20000 2924 20052
rect 3056 19864 3108 19916
rect 7472 20000 7524 20052
rect 8116 20000 8168 20052
rect 3792 19796 3844 19848
rect 3884 19796 3936 19848
rect 4804 19907 4856 19916
rect 4804 19873 4813 19907
rect 4813 19873 4847 19907
rect 4847 19873 4856 19907
rect 4804 19864 4856 19873
rect 5908 19796 5960 19848
rect 7932 19932 7984 19984
rect 10232 20000 10284 20052
rect 11612 20043 11664 20052
rect 11612 20009 11621 20043
rect 11621 20009 11655 20043
rect 11655 20009 11664 20043
rect 11612 20000 11664 20009
rect 14004 20000 14056 20052
rect 14096 20000 14148 20052
rect 1768 19703 1820 19712
rect 1768 19669 1777 19703
rect 1777 19669 1811 19703
rect 1811 19669 1820 19703
rect 1768 19660 1820 19669
rect 2964 19660 3016 19712
rect 3976 19660 4028 19712
rect 4620 19728 4672 19780
rect 5080 19660 5132 19712
rect 5172 19703 5224 19712
rect 5172 19669 5181 19703
rect 5181 19669 5215 19703
rect 5215 19669 5224 19703
rect 5172 19660 5224 19669
rect 6552 19839 6604 19848
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 6644 19839 6696 19848
rect 6644 19805 6653 19839
rect 6653 19805 6687 19839
rect 6687 19805 6696 19839
rect 6644 19796 6696 19805
rect 8392 19796 8444 19848
rect 6920 19771 6972 19780
rect 6920 19737 6929 19771
rect 6929 19737 6963 19771
rect 6963 19737 6972 19771
rect 6920 19728 6972 19737
rect 8300 19728 8352 19780
rect 7564 19660 7616 19712
rect 9312 19796 9364 19848
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 9588 19839 9640 19848
rect 9588 19805 9597 19839
rect 9597 19805 9631 19839
rect 9631 19805 9640 19839
rect 9588 19796 9640 19805
rect 9680 19796 9732 19848
rect 11796 19932 11848 19984
rect 12900 19975 12952 19984
rect 12900 19941 12909 19975
rect 12909 19941 12943 19975
rect 12943 19941 12952 19975
rect 12900 19932 12952 19941
rect 13452 19932 13504 19984
rect 14372 19932 14424 19984
rect 16120 20000 16172 20052
rect 15844 19975 15896 19984
rect 15844 19941 15853 19975
rect 15853 19941 15887 19975
rect 15887 19941 15896 19975
rect 15844 19932 15896 19941
rect 16856 20043 16908 20052
rect 16856 20009 16865 20043
rect 16865 20009 16899 20043
rect 16899 20009 16908 20043
rect 16856 20000 16908 20009
rect 17684 20000 17736 20052
rect 17960 20000 18012 20052
rect 18236 20000 18288 20052
rect 18696 20000 18748 20052
rect 20812 20000 20864 20052
rect 22192 20000 22244 20052
rect 22928 20000 22980 20052
rect 23388 20000 23440 20052
rect 24124 20000 24176 20052
rect 26332 20043 26384 20052
rect 26332 20009 26341 20043
rect 26341 20009 26375 20043
rect 26375 20009 26384 20043
rect 26332 20000 26384 20009
rect 26424 20043 26476 20052
rect 26424 20009 26433 20043
rect 26433 20009 26467 20043
rect 26467 20009 26476 20043
rect 26424 20000 26476 20009
rect 28632 20000 28684 20052
rect 28816 20000 28868 20052
rect 28908 20000 28960 20052
rect 29736 20000 29788 20052
rect 16580 19932 16632 19984
rect 17776 19932 17828 19984
rect 9956 19796 10008 19848
rect 10140 19839 10192 19848
rect 10140 19805 10149 19839
rect 10149 19805 10183 19839
rect 10183 19805 10192 19839
rect 10140 19796 10192 19805
rect 12072 19796 12124 19848
rect 12532 19796 12584 19848
rect 13728 19796 13780 19848
rect 14004 19796 14056 19848
rect 8944 19660 8996 19712
rect 9772 19660 9824 19712
rect 11428 19703 11480 19712
rect 11428 19669 11437 19703
rect 11437 19669 11471 19703
rect 11471 19669 11480 19703
rect 11428 19660 11480 19669
rect 11796 19660 11848 19712
rect 13360 19660 13412 19712
rect 13452 19703 13504 19712
rect 13452 19669 13461 19703
rect 13461 19669 13495 19703
rect 13495 19669 13504 19703
rect 13452 19660 13504 19669
rect 13636 19771 13688 19780
rect 13636 19737 13645 19771
rect 13645 19737 13679 19771
rect 13679 19737 13688 19771
rect 14740 19864 14792 19916
rect 15476 19796 15528 19848
rect 15660 19839 15712 19848
rect 15660 19805 15669 19839
rect 15669 19805 15703 19839
rect 15703 19805 15712 19839
rect 15660 19796 15712 19805
rect 16212 19796 16264 19848
rect 16304 19839 16356 19848
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 16396 19839 16448 19848
rect 16396 19805 16405 19839
rect 16405 19805 16439 19839
rect 16439 19805 16448 19839
rect 16396 19796 16448 19805
rect 16856 19796 16908 19848
rect 20076 19864 20128 19916
rect 20996 19864 21048 19916
rect 23848 19907 23900 19916
rect 23848 19873 23857 19907
rect 23857 19873 23891 19907
rect 23891 19873 23900 19907
rect 23848 19864 23900 19873
rect 23940 19864 23992 19916
rect 17408 19839 17460 19848
rect 17408 19805 17417 19839
rect 17417 19805 17451 19839
rect 17451 19805 17460 19839
rect 17408 19796 17460 19805
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 13636 19728 13688 19737
rect 16580 19728 16632 19780
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 18696 19796 18748 19805
rect 19064 19796 19116 19848
rect 19892 19839 19944 19848
rect 19892 19805 19901 19839
rect 19901 19805 19935 19839
rect 19935 19805 19944 19839
rect 19892 19796 19944 19805
rect 19984 19839 20036 19848
rect 19984 19805 19993 19839
rect 19993 19805 20027 19839
rect 20027 19805 20036 19839
rect 19984 19796 20036 19805
rect 18236 19728 18288 19780
rect 19248 19728 19300 19780
rect 20352 19796 20404 19848
rect 20536 19839 20588 19848
rect 20536 19805 20545 19839
rect 20545 19805 20579 19839
rect 20579 19805 20588 19839
rect 20536 19796 20588 19805
rect 14004 19660 14056 19712
rect 17960 19660 18012 19712
rect 18144 19660 18196 19712
rect 20812 19728 20864 19780
rect 18880 19660 18932 19712
rect 20168 19660 20220 19712
rect 20628 19660 20680 19712
rect 22652 19796 22704 19848
rect 23296 19796 23348 19848
rect 23388 19796 23440 19848
rect 23572 19796 23624 19848
rect 26332 19864 26384 19916
rect 22836 19771 22888 19780
rect 22836 19737 22845 19771
rect 22845 19737 22879 19771
rect 22879 19737 22888 19771
rect 22836 19728 22888 19737
rect 23480 19703 23532 19712
rect 23480 19669 23489 19703
rect 23489 19669 23523 19703
rect 23523 19669 23532 19703
rect 23480 19660 23532 19669
rect 23572 19660 23624 19712
rect 24492 19796 24544 19848
rect 24676 19796 24728 19848
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 24860 19728 24912 19780
rect 25136 19796 25188 19848
rect 25504 19796 25556 19848
rect 25872 19796 25924 19848
rect 25228 19771 25280 19780
rect 25228 19737 25237 19771
rect 25237 19737 25271 19771
rect 25271 19737 25280 19771
rect 25228 19728 25280 19737
rect 25320 19771 25372 19780
rect 25320 19737 25329 19771
rect 25329 19737 25363 19771
rect 25363 19737 25372 19771
rect 25320 19728 25372 19737
rect 26700 19839 26752 19848
rect 26700 19805 26709 19839
rect 26709 19805 26743 19839
rect 26743 19805 26752 19839
rect 26700 19796 26752 19805
rect 27160 19796 27212 19848
rect 27252 19796 27304 19848
rect 28724 19864 28776 19916
rect 29552 19864 29604 19916
rect 26792 19771 26844 19780
rect 26792 19737 26801 19771
rect 26801 19737 26835 19771
rect 26835 19737 26844 19771
rect 26792 19728 26844 19737
rect 28540 19771 28592 19780
rect 28540 19737 28549 19771
rect 28549 19737 28583 19771
rect 28583 19737 28592 19771
rect 28540 19728 28592 19737
rect 29644 19796 29696 19848
rect 29828 19839 29880 19848
rect 29828 19805 29837 19839
rect 29837 19805 29871 19839
rect 29871 19805 29880 19839
rect 29828 19796 29880 19805
rect 30656 20000 30708 20052
rect 32036 20000 32088 20052
rect 34704 20000 34756 20052
rect 35164 20000 35216 20052
rect 35716 20000 35768 20052
rect 35808 20000 35860 20052
rect 29368 19728 29420 19780
rect 30196 19728 30248 19780
rect 30748 19864 30800 19916
rect 31208 19907 31260 19916
rect 31208 19873 31217 19907
rect 31217 19873 31251 19907
rect 31251 19873 31260 19907
rect 31208 19864 31260 19873
rect 31576 19796 31628 19848
rect 34612 19932 34664 19984
rect 32956 19864 33008 19916
rect 33140 19864 33192 19916
rect 35164 19839 35216 19848
rect 35164 19805 35173 19839
rect 35173 19805 35207 19839
rect 35207 19805 35216 19839
rect 35164 19796 35216 19805
rect 35440 19839 35492 19848
rect 35440 19805 35449 19839
rect 35449 19805 35483 19839
rect 35483 19805 35492 19839
rect 35440 19796 35492 19805
rect 35624 19864 35676 19916
rect 28954 19660 29006 19712
rect 29184 19660 29236 19712
rect 29552 19703 29604 19712
rect 29552 19669 29561 19703
rect 29561 19669 29595 19703
rect 29595 19669 29604 19703
rect 29552 19660 29604 19669
rect 34796 19660 34848 19712
rect 35900 19703 35952 19712
rect 35900 19669 35909 19703
rect 35909 19669 35943 19703
rect 35943 19669 35952 19703
rect 35900 19660 35952 19669
rect 36176 19660 36228 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1400 19456 1452 19508
rect 1768 19388 1820 19440
rect 2964 19388 3016 19440
rect 3608 19320 3660 19372
rect 3884 19431 3936 19440
rect 3884 19397 3893 19431
rect 3893 19397 3927 19431
rect 3927 19397 3936 19431
rect 3884 19388 3936 19397
rect 5080 19456 5132 19508
rect 5908 19499 5960 19508
rect 5908 19465 5917 19499
rect 5917 19465 5951 19499
rect 5951 19465 5960 19499
rect 5908 19456 5960 19465
rect 6552 19456 6604 19508
rect 6920 19456 6972 19508
rect 7196 19456 7248 19508
rect 8208 19456 8260 19508
rect 9588 19456 9640 19508
rect 3148 19227 3200 19236
rect 3148 19193 3157 19227
rect 3157 19193 3191 19227
rect 3191 19193 3200 19227
rect 3148 19184 3200 19193
rect 5448 19320 5500 19372
rect 8944 19431 8996 19440
rect 8944 19397 8953 19431
rect 8953 19397 8987 19431
rect 8987 19397 8996 19431
rect 8944 19388 8996 19397
rect 9036 19431 9088 19440
rect 9036 19397 9045 19431
rect 9045 19397 9079 19431
rect 9079 19397 9088 19431
rect 9036 19388 9088 19397
rect 3976 19252 4028 19304
rect 4804 19252 4856 19304
rect 8208 19320 8260 19372
rect 8760 19363 8812 19372
rect 8760 19329 8769 19363
rect 8769 19329 8803 19363
rect 8803 19329 8812 19363
rect 8760 19320 8812 19329
rect 9496 19320 9548 19372
rect 11796 19456 11848 19508
rect 9956 19320 10008 19372
rect 11060 19320 11112 19372
rect 8300 19295 8352 19304
rect 8300 19261 8309 19295
rect 8309 19261 8343 19295
rect 8343 19261 8352 19295
rect 8300 19252 8352 19261
rect 9312 19252 9364 19304
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 13176 19499 13228 19508
rect 13176 19465 13185 19499
rect 13185 19465 13219 19499
rect 13219 19465 13228 19499
rect 13176 19456 13228 19465
rect 12164 19388 12216 19440
rect 13728 19388 13780 19440
rect 12256 19363 12308 19372
rect 12256 19329 12265 19363
rect 12265 19329 12299 19363
rect 12299 19329 12308 19363
rect 12256 19320 12308 19329
rect 12532 19363 12584 19372
rect 12532 19329 12541 19363
rect 12541 19329 12575 19363
rect 12575 19329 12584 19363
rect 12532 19320 12584 19329
rect 9220 19184 9272 19236
rect 11796 19295 11848 19304
rect 11796 19261 11805 19295
rect 11805 19261 11839 19295
rect 11839 19261 11848 19295
rect 11796 19252 11848 19261
rect 12072 19252 12124 19304
rect 13360 19363 13412 19372
rect 13360 19329 13369 19363
rect 13369 19329 13403 19363
rect 13403 19329 13412 19363
rect 13360 19320 13412 19329
rect 14280 19363 14332 19372
rect 14280 19329 14289 19363
rect 14289 19329 14323 19363
rect 14323 19329 14332 19363
rect 14280 19320 14332 19329
rect 15660 19456 15712 19508
rect 15844 19456 15896 19508
rect 16212 19456 16264 19508
rect 14740 19363 14792 19372
rect 14740 19329 14749 19363
rect 14749 19329 14783 19363
rect 14783 19329 14792 19363
rect 14740 19320 14792 19329
rect 16304 19388 16356 19440
rect 18144 19456 18196 19508
rect 19524 19456 19576 19508
rect 19984 19456 20036 19508
rect 22100 19456 22152 19508
rect 17408 19320 17460 19372
rect 19248 19388 19300 19440
rect 19340 19320 19392 19372
rect 19616 19320 19668 19372
rect 21916 19388 21968 19440
rect 19984 19320 20036 19372
rect 20536 19320 20588 19372
rect 13912 19252 13964 19304
rect 11336 19159 11388 19168
rect 11336 19125 11345 19159
rect 11345 19125 11379 19159
rect 11379 19125 11388 19159
rect 11336 19116 11388 19125
rect 12164 19184 12216 19236
rect 14648 19227 14700 19236
rect 14648 19193 14657 19227
rect 14657 19193 14691 19227
rect 14691 19193 14700 19227
rect 14648 19184 14700 19193
rect 16764 19227 16816 19236
rect 16764 19193 16773 19227
rect 16773 19193 16807 19227
rect 16807 19193 16816 19227
rect 16764 19184 16816 19193
rect 17776 19252 17828 19304
rect 20168 19252 20220 19304
rect 22376 19388 22428 19440
rect 22836 19456 22888 19508
rect 23848 19499 23900 19508
rect 23848 19465 23857 19499
rect 23857 19465 23891 19499
rect 23891 19465 23900 19499
rect 23848 19456 23900 19465
rect 23940 19456 23992 19508
rect 24768 19456 24820 19508
rect 25872 19456 25924 19508
rect 27160 19456 27212 19508
rect 28080 19456 28132 19508
rect 28724 19456 28776 19508
rect 29184 19456 29236 19508
rect 29552 19456 29604 19508
rect 29736 19456 29788 19508
rect 29828 19456 29880 19508
rect 30380 19456 30432 19508
rect 32956 19456 33008 19508
rect 23480 19388 23532 19440
rect 22560 19320 22612 19372
rect 23112 19320 23164 19372
rect 23388 19320 23440 19372
rect 24492 19388 24544 19440
rect 27068 19388 27120 19440
rect 27436 19431 27488 19440
rect 27436 19397 27445 19431
rect 27445 19397 27479 19431
rect 27479 19397 27488 19431
rect 27436 19388 27488 19397
rect 27528 19431 27580 19440
rect 27528 19397 27537 19431
rect 27537 19397 27571 19431
rect 27571 19397 27580 19431
rect 27528 19388 27580 19397
rect 27988 19388 28040 19440
rect 27252 19363 27304 19372
rect 27252 19329 27281 19363
rect 27281 19329 27304 19363
rect 27252 19320 27304 19329
rect 24308 19295 24360 19304
rect 24308 19261 24317 19295
rect 24317 19261 24351 19295
rect 24351 19261 24360 19295
rect 27620 19363 27672 19372
rect 27620 19329 27629 19363
rect 27629 19329 27663 19363
rect 27663 19329 27672 19363
rect 27620 19320 27672 19329
rect 27804 19320 27856 19372
rect 28080 19363 28132 19372
rect 28080 19329 28089 19363
rect 28089 19329 28123 19363
rect 28123 19329 28132 19363
rect 28080 19320 28132 19329
rect 28264 19363 28316 19372
rect 28264 19329 28273 19363
rect 28273 19329 28307 19363
rect 28307 19329 28316 19363
rect 28264 19320 28316 19329
rect 28540 19320 28592 19372
rect 29368 19363 29420 19372
rect 29368 19329 29377 19363
rect 29377 19329 29411 19363
rect 29411 19329 29420 19363
rect 29368 19320 29420 19329
rect 29552 19320 29604 19372
rect 33140 19363 33192 19372
rect 33140 19329 33149 19363
rect 33149 19329 33183 19363
rect 33183 19329 33192 19363
rect 33140 19320 33192 19329
rect 24308 19252 24360 19261
rect 28172 19252 28224 19304
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 12900 19116 12952 19125
rect 17224 19116 17276 19168
rect 22100 19116 22152 19168
rect 25688 19184 25740 19236
rect 24124 19116 24176 19168
rect 26792 19116 26844 19168
rect 29644 19159 29696 19168
rect 29644 19125 29653 19159
rect 29653 19125 29687 19159
rect 29687 19125 29696 19159
rect 29644 19116 29696 19125
rect 33140 19159 33192 19168
rect 33140 19125 33149 19159
rect 33149 19125 33183 19159
rect 33183 19125 33192 19159
rect 34152 19363 34204 19372
rect 34152 19329 34161 19363
rect 34161 19329 34195 19363
rect 34195 19329 34204 19363
rect 34152 19320 34204 19329
rect 34796 19456 34848 19508
rect 35900 19499 35952 19508
rect 35900 19465 35909 19499
rect 35909 19465 35943 19499
rect 35943 19465 35952 19499
rect 35900 19456 35952 19465
rect 34796 19295 34848 19304
rect 34796 19261 34805 19295
rect 34805 19261 34839 19295
rect 34839 19261 34848 19295
rect 34796 19252 34848 19261
rect 34428 19184 34480 19236
rect 33140 19116 33192 19125
rect 35992 19116 36044 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4804 18912 4856 18964
rect 17224 18912 17276 18964
rect 18052 18912 18104 18964
rect 18972 18912 19024 18964
rect 4068 18776 4120 18828
rect 5908 18776 5960 18828
rect 13912 18844 13964 18896
rect 10876 18819 10928 18828
rect 10876 18785 10885 18819
rect 10885 18785 10919 18819
rect 10919 18785 10928 18819
rect 10876 18776 10928 18785
rect 11428 18776 11480 18828
rect 5172 18708 5224 18760
rect 6000 18751 6052 18760
rect 6000 18717 6009 18751
rect 6009 18717 6043 18751
rect 6043 18717 6052 18751
rect 6000 18708 6052 18717
rect 11888 18751 11940 18760
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 11888 18708 11940 18717
rect 12072 18708 12124 18760
rect 940 18640 992 18692
rect 1768 18683 1820 18692
rect 1768 18649 1777 18683
rect 1777 18649 1811 18683
rect 1811 18649 1820 18683
rect 1768 18640 1820 18649
rect 3148 18640 3200 18692
rect 5632 18683 5684 18692
rect 5632 18649 5641 18683
rect 5641 18649 5675 18683
rect 5675 18649 5684 18683
rect 5632 18640 5684 18649
rect 5816 18640 5868 18692
rect 9220 18640 9272 18692
rect 1952 18572 2004 18624
rect 4252 18572 4304 18624
rect 6552 18572 6604 18624
rect 6736 18572 6788 18624
rect 10048 18572 10100 18624
rect 10324 18615 10376 18624
rect 10324 18581 10333 18615
rect 10333 18581 10367 18615
rect 10367 18581 10376 18615
rect 10324 18572 10376 18581
rect 11336 18572 11388 18624
rect 12348 18708 12400 18760
rect 18604 18844 18656 18896
rect 19432 18912 19484 18964
rect 19984 18912 20036 18964
rect 20168 18912 20220 18964
rect 20720 18912 20772 18964
rect 20904 18912 20956 18964
rect 21088 18912 21140 18964
rect 22652 18912 22704 18964
rect 23204 18912 23256 18964
rect 26792 18912 26844 18964
rect 32864 18912 32916 18964
rect 34428 18912 34480 18964
rect 19340 18819 19392 18828
rect 19340 18785 19349 18819
rect 19349 18785 19383 18819
rect 19383 18785 19392 18819
rect 19340 18776 19392 18785
rect 16764 18708 16816 18760
rect 17684 18751 17736 18760
rect 17684 18717 17693 18751
rect 17693 18717 17727 18751
rect 17727 18717 17736 18751
rect 17684 18708 17736 18717
rect 12532 18640 12584 18692
rect 13360 18640 13412 18692
rect 17132 18640 17184 18692
rect 18052 18751 18104 18760
rect 18052 18717 18061 18751
rect 18061 18717 18095 18751
rect 18095 18717 18104 18751
rect 18052 18708 18104 18717
rect 18420 18708 18472 18760
rect 18696 18640 18748 18692
rect 19248 18751 19300 18760
rect 19248 18717 19257 18751
rect 19257 18717 19291 18751
rect 19291 18717 19300 18751
rect 19248 18708 19300 18717
rect 19524 18751 19576 18760
rect 19524 18717 19533 18751
rect 19533 18717 19567 18751
rect 19567 18717 19576 18751
rect 19524 18708 19576 18717
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 19984 18819 20036 18828
rect 19984 18785 19993 18819
rect 19993 18785 20027 18819
rect 20027 18785 20036 18819
rect 19984 18776 20036 18785
rect 14188 18615 14240 18624
rect 14188 18581 14197 18615
rect 14197 18581 14231 18615
rect 14231 18581 14240 18615
rect 14188 18572 14240 18581
rect 15476 18572 15528 18624
rect 15752 18572 15804 18624
rect 18052 18615 18104 18624
rect 18052 18581 18061 18615
rect 18061 18581 18095 18615
rect 18095 18581 18104 18615
rect 18052 18572 18104 18581
rect 18788 18572 18840 18624
rect 18880 18572 18932 18624
rect 20628 18708 20680 18760
rect 25872 18844 25924 18896
rect 27436 18844 27488 18896
rect 23480 18776 23532 18828
rect 21640 18751 21692 18760
rect 21640 18717 21649 18751
rect 21649 18717 21683 18751
rect 21683 18717 21692 18751
rect 21640 18708 21692 18717
rect 22376 18751 22428 18760
rect 22376 18717 22385 18751
rect 22385 18717 22419 18751
rect 22419 18717 22428 18751
rect 22376 18708 22428 18717
rect 21180 18683 21232 18692
rect 21180 18649 21189 18683
rect 21189 18649 21223 18683
rect 21223 18649 21232 18683
rect 21180 18640 21232 18649
rect 31300 18708 31352 18760
rect 31392 18751 31444 18760
rect 31392 18717 31401 18751
rect 31401 18717 31435 18751
rect 31435 18717 31444 18751
rect 31392 18708 31444 18717
rect 33140 18776 33192 18828
rect 32680 18751 32732 18760
rect 32680 18717 32689 18751
rect 32689 18717 32723 18751
rect 32723 18717 32732 18751
rect 32680 18708 32732 18717
rect 32772 18751 32824 18760
rect 32772 18717 32781 18751
rect 32781 18717 32815 18751
rect 32815 18717 32824 18751
rect 32772 18708 32824 18717
rect 32956 18708 33008 18760
rect 33968 18708 34020 18760
rect 35440 18776 35492 18828
rect 36728 18819 36780 18828
rect 36728 18785 36737 18819
rect 36737 18785 36771 18819
rect 36771 18785 36780 18819
rect 36728 18776 36780 18785
rect 36820 18640 36872 18692
rect 20996 18615 21048 18624
rect 20996 18581 21023 18615
rect 21023 18581 21048 18615
rect 20996 18572 21048 18581
rect 22192 18615 22244 18624
rect 22192 18581 22201 18615
rect 22201 18581 22235 18615
rect 22235 18581 22244 18615
rect 22192 18572 22244 18581
rect 25596 18572 25648 18624
rect 26056 18572 26108 18624
rect 28448 18572 28500 18624
rect 30748 18572 30800 18624
rect 31024 18572 31076 18624
rect 31208 18615 31260 18624
rect 31208 18581 31217 18615
rect 31217 18581 31251 18615
rect 31251 18581 31260 18615
rect 31208 18572 31260 18581
rect 32312 18572 32364 18624
rect 32956 18572 33008 18624
rect 33140 18572 33192 18624
rect 34796 18615 34848 18624
rect 34796 18581 34811 18615
rect 34811 18581 34845 18615
rect 34845 18581 34848 18615
rect 34796 18572 34848 18581
rect 34980 18572 35032 18624
rect 35164 18572 35216 18624
rect 37096 18615 37148 18624
rect 37096 18581 37105 18615
rect 37105 18581 37139 18615
rect 37139 18581 37148 18615
rect 37096 18572 37148 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4252 18368 4304 18420
rect 8300 18300 8352 18352
rect 10232 18300 10284 18352
rect 10784 18300 10836 18352
rect 13820 18368 13872 18420
rect 13912 18411 13964 18420
rect 13912 18377 13921 18411
rect 13921 18377 13955 18411
rect 13955 18377 13964 18411
rect 13912 18368 13964 18377
rect 14188 18368 14240 18420
rect 15384 18411 15436 18420
rect 15384 18377 15393 18411
rect 15393 18377 15427 18411
rect 15427 18377 15436 18411
rect 15384 18368 15436 18377
rect 19340 18368 19392 18420
rect 11336 18300 11388 18352
rect 12256 18300 12308 18352
rect 1676 18207 1728 18216
rect 1676 18173 1685 18207
rect 1685 18173 1719 18207
rect 1719 18173 1728 18207
rect 1676 18164 1728 18173
rect 6736 18232 6788 18284
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 12532 18275 12584 18284
rect 12532 18241 12541 18275
rect 12541 18241 12575 18275
rect 12575 18241 12584 18275
rect 12532 18232 12584 18241
rect 12808 18232 12860 18284
rect 14004 18232 14056 18284
rect 14188 18232 14240 18284
rect 16856 18300 16908 18352
rect 16396 18232 16448 18284
rect 17040 18232 17092 18284
rect 17592 18300 17644 18352
rect 18420 18300 18472 18352
rect 18236 18232 18288 18284
rect 19064 18300 19116 18352
rect 22100 18368 22152 18420
rect 19984 18300 20036 18352
rect 4068 18164 4120 18216
rect 5908 18207 5960 18216
rect 5908 18173 5917 18207
rect 5917 18173 5951 18207
rect 5951 18173 5960 18207
rect 5908 18164 5960 18173
rect 3700 18096 3752 18148
rect 6644 18164 6696 18216
rect 2044 18071 2096 18080
rect 2044 18037 2053 18071
rect 2053 18037 2087 18071
rect 2087 18037 2096 18071
rect 2044 18028 2096 18037
rect 2504 18071 2556 18080
rect 2504 18037 2513 18071
rect 2513 18037 2547 18071
rect 2547 18037 2556 18071
rect 2504 18028 2556 18037
rect 2964 18028 3016 18080
rect 3516 18028 3568 18080
rect 6184 18028 6236 18080
rect 7932 18164 7984 18216
rect 9220 18164 9272 18216
rect 10784 18096 10836 18148
rect 11152 18096 11204 18148
rect 12072 18164 12124 18216
rect 12716 18164 12768 18216
rect 13912 18164 13964 18216
rect 14740 18207 14792 18216
rect 14740 18173 14749 18207
rect 14749 18173 14783 18207
rect 14783 18173 14792 18207
rect 14740 18164 14792 18173
rect 15568 18207 15620 18216
rect 15568 18173 15577 18207
rect 15577 18173 15611 18207
rect 15611 18173 15620 18207
rect 15568 18164 15620 18173
rect 15476 18096 15528 18148
rect 15936 18164 15988 18216
rect 18972 18232 19024 18284
rect 19432 18164 19484 18216
rect 19616 18275 19668 18284
rect 19616 18241 19626 18275
rect 19626 18241 19660 18275
rect 19660 18241 19668 18275
rect 19616 18232 19668 18241
rect 20444 18232 20496 18284
rect 22376 18232 22428 18284
rect 22652 18300 22704 18352
rect 29460 18300 29512 18352
rect 22560 18232 22612 18284
rect 23940 18232 23992 18284
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 25136 18232 25188 18284
rect 23664 18164 23716 18216
rect 25412 18275 25464 18284
rect 25412 18241 25421 18275
rect 25421 18241 25455 18275
rect 25455 18241 25464 18275
rect 25412 18232 25464 18241
rect 26056 18232 26108 18284
rect 27988 18275 28040 18284
rect 27988 18241 27997 18275
rect 27997 18241 28031 18275
rect 28031 18241 28040 18275
rect 27988 18232 28040 18241
rect 28172 18275 28224 18284
rect 28172 18241 28181 18275
rect 28181 18241 28215 18275
rect 28215 18241 28224 18275
rect 28172 18232 28224 18241
rect 30380 18300 30432 18352
rect 31208 18368 31260 18420
rect 25780 18207 25832 18216
rect 25780 18173 25789 18207
rect 25789 18173 25823 18207
rect 25823 18173 25832 18207
rect 25780 18164 25832 18173
rect 28632 18164 28684 18216
rect 8852 18028 8904 18080
rect 9128 18028 9180 18080
rect 14280 18028 14332 18080
rect 14648 18028 14700 18080
rect 15384 18028 15436 18080
rect 16948 18028 17000 18080
rect 17960 18028 18012 18080
rect 18512 18028 18564 18080
rect 18880 18028 18932 18080
rect 19248 18028 19300 18080
rect 19616 18028 19668 18080
rect 24676 18096 24728 18148
rect 25688 18096 25740 18148
rect 26240 18139 26292 18148
rect 26240 18105 26249 18139
rect 26249 18105 26283 18139
rect 26283 18105 26292 18139
rect 26240 18096 26292 18105
rect 28908 18096 28960 18148
rect 29920 18164 29972 18216
rect 30840 18232 30892 18284
rect 31300 18300 31352 18352
rect 32680 18368 32732 18420
rect 34152 18368 34204 18420
rect 34796 18368 34848 18420
rect 37096 18368 37148 18420
rect 31024 18275 31076 18284
rect 31024 18241 31033 18275
rect 31033 18241 31067 18275
rect 31067 18241 31076 18275
rect 31024 18232 31076 18241
rect 32036 18232 32088 18284
rect 33140 18343 33192 18352
rect 33140 18309 33149 18343
rect 33149 18309 33183 18343
rect 33183 18309 33192 18343
rect 33140 18300 33192 18309
rect 32680 18232 32732 18284
rect 31576 18164 31628 18216
rect 32496 18207 32548 18216
rect 32496 18173 32505 18207
rect 32505 18173 32539 18207
rect 32539 18173 32548 18207
rect 32496 18164 32548 18173
rect 32588 18207 32640 18216
rect 32588 18173 32597 18207
rect 32597 18173 32631 18207
rect 32631 18173 32640 18207
rect 32588 18164 32640 18173
rect 32128 18096 32180 18148
rect 32772 18096 32824 18148
rect 26516 18028 26568 18080
rect 27896 18028 27948 18080
rect 29552 18071 29604 18080
rect 29552 18037 29561 18071
rect 29561 18037 29595 18071
rect 29595 18037 29604 18071
rect 29552 18028 29604 18037
rect 29920 18028 29972 18080
rect 31760 18028 31812 18080
rect 34980 18275 35032 18284
rect 34980 18241 34989 18275
rect 34989 18241 35023 18275
rect 35023 18241 35032 18275
rect 34980 18232 35032 18241
rect 35624 18300 35676 18352
rect 35164 18275 35216 18284
rect 35164 18241 35173 18275
rect 35173 18241 35207 18275
rect 35207 18241 35216 18275
rect 35164 18232 35216 18241
rect 37188 18300 37240 18352
rect 33968 18028 34020 18080
rect 37556 18028 37608 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 38384 17960 38436 18012
rect 1768 17824 1820 17876
rect 2136 17824 2188 17876
rect 1676 17688 1728 17740
rect 1952 17620 2004 17672
rect 2044 17620 2096 17672
rect 5632 17824 5684 17876
rect 6920 17824 6972 17876
rect 7748 17824 7800 17876
rect 7932 17824 7984 17876
rect 8300 17756 8352 17808
rect 3516 17688 3568 17740
rect 3976 17731 4028 17740
rect 3976 17697 3985 17731
rect 3985 17697 4019 17731
rect 4019 17697 4028 17731
rect 3976 17688 4028 17697
rect 5448 17688 5500 17740
rect 9864 17824 9916 17876
rect 11704 17824 11756 17876
rect 12440 17867 12492 17876
rect 12440 17833 12449 17867
rect 12449 17833 12483 17867
rect 12483 17833 12492 17867
rect 12440 17824 12492 17833
rect 12532 17824 12584 17876
rect 13084 17824 13136 17876
rect 14740 17824 14792 17876
rect 15200 17824 15252 17876
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 3700 17620 3752 17672
rect 4252 17595 4304 17604
rect 4252 17561 4261 17595
rect 4261 17561 4295 17595
rect 4295 17561 4304 17595
rect 4252 17552 4304 17561
rect 9128 17688 9180 17740
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 11152 17688 11204 17740
rect 11612 17688 11664 17740
rect 11980 17731 12032 17740
rect 11980 17697 11989 17731
rect 11989 17697 12023 17731
rect 12023 17697 12032 17731
rect 11980 17688 12032 17697
rect 6368 17595 6420 17604
rect 6368 17561 6377 17595
rect 6377 17561 6411 17595
rect 6411 17561 6420 17595
rect 6368 17552 6420 17561
rect 6920 17552 6972 17604
rect 5724 17527 5776 17536
rect 5724 17493 5733 17527
rect 5733 17493 5767 17527
rect 5767 17493 5776 17527
rect 5724 17484 5776 17493
rect 6184 17484 6236 17536
rect 7196 17484 7248 17536
rect 7380 17484 7432 17536
rect 10324 17620 10376 17672
rect 10508 17620 10560 17672
rect 10600 17620 10652 17672
rect 11060 17663 11112 17672
rect 11060 17629 11069 17663
rect 11069 17629 11103 17663
rect 11103 17629 11112 17663
rect 11060 17620 11112 17629
rect 11888 17620 11940 17672
rect 12348 17620 12400 17672
rect 9588 17484 9640 17536
rect 12532 17731 12584 17740
rect 12532 17697 12541 17731
rect 12541 17697 12575 17731
rect 12575 17697 12584 17731
rect 12532 17688 12584 17697
rect 13360 17688 13412 17740
rect 14648 17731 14700 17740
rect 14648 17697 14657 17731
rect 14657 17697 14691 17731
rect 14691 17697 14700 17731
rect 14648 17688 14700 17697
rect 15108 17688 15160 17740
rect 12808 17552 12860 17604
rect 14188 17620 14240 17672
rect 12164 17484 12216 17536
rect 12256 17527 12308 17536
rect 12256 17493 12265 17527
rect 12265 17493 12299 17527
rect 12299 17493 12308 17527
rect 12256 17484 12308 17493
rect 12348 17484 12400 17536
rect 13084 17484 13136 17536
rect 13636 17527 13688 17536
rect 13636 17493 13645 17527
rect 13645 17493 13679 17527
rect 13679 17493 13688 17527
rect 13636 17484 13688 17493
rect 14004 17484 14056 17536
rect 14464 17620 14516 17672
rect 15752 17688 15804 17740
rect 20812 17824 20864 17876
rect 21640 17824 21692 17876
rect 22744 17824 22796 17876
rect 23296 17824 23348 17876
rect 26884 17824 26936 17876
rect 17224 17756 17276 17808
rect 23664 17756 23716 17808
rect 14372 17552 14424 17604
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 16120 17620 16172 17672
rect 16580 17688 16632 17740
rect 15384 17552 15436 17604
rect 15752 17552 15804 17604
rect 16764 17620 16816 17672
rect 16948 17620 17000 17672
rect 17684 17663 17736 17672
rect 17684 17629 17693 17663
rect 17693 17629 17727 17663
rect 17727 17629 17736 17663
rect 17684 17620 17736 17629
rect 17040 17552 17092 17604
rect 17776 17552 17828 17604
rect 18052 17663 18104 17672
rect 18052 17629 18061 17663
rect 18061 17629 18095 17663
rect 18095 17629 18104 17663
rect 18052 17620 18104 17629
rect 18144 17663 18196 17672
rect 18144 17629 18153 17663
rect 18153 17629 18187 17663
rect 18187 17629 18196 17663
rect 18144 17620 18196 17629
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 18604 17620 18656 17672
rect 18696 17620 18748 17672
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 19340 17620 19392 17672
rect 19432 17620 19484 17672
rect 19984 17620 20036 17672
rect 20168 17620 20220 17672
rect 21180 17620 21232 17672
rect 22100 17620 22152 17672
rect 22284 17663 22336 17672
rect 22284 17629 22293 17663
rect 22293 17629 22327 17663
rect 22327 17629 22336 17663
rect 22284 17620 22336 17629
rect 23480 17731 23532 17740
rect 23480 17697 23489 17731
rect 23489 17697 23523 17731
rect 23523 17697 23532 17731
rect 23480 17688 23532 17697
rect 24676 17731 24728 17740
rect 24676 17697 24685 17731
rect 24685 17697 24719 17731
rect 24719 17697 24728 17731
rect 24676 17688 24728 17697
rect 17316 17484 17368 17536
rect 20628 17552 20680 17604
rect 24032 17620 24084 17672
rect 24768 17620 24820 17672
rect 26240 17756 26292 17808
rect 27988 17824 28040 17876
rect 31208 17824 31260 17876
rect 31392 17824 31444 17876
rect 32496 17824 32548 17876
rect 27712 17731 27764 17740
rect 27712 17697 27721 17731
rect 27721 17697 27755 17731
rect 27755 17697 27764 17731
rect 27712 17688 27764 17697
rect 29828 17756 29880 17808
rect 28264 17688 28316 17740
rect 27804 17620 27856 17672
rect 27896 17663 27948 17672
rect 27896 17629 27905 17663
rect 27905 17629 27939 17663
rect 27939 17629 27948 17663
rect 27896 17620 27948 17629
rect 27988 17620 28040 17672
rect 28356 17663 28408 17672
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 27344 17552 27396 17604
rect 28172 17552 28224 17604
rect 28632 17620 28684 17672
rect 29736 17663 29788 17672
rect 29736 17629 29745 17663
rect 29745 17629 29779 17663
rect 29779 17629 29788 17663
rect 29736 17620 29788 17629
rect 30104 17620 30156 17672
rect 30288 17756 30340 17808
rect 30288 17663 30340 17672
rect 30288 17629 30297 17663
rect 30297 17629 30331 17663
rect 30331 17629 30340 17663
rect 30288 17620 30340 17629
rect 32588 17756 32640 17808
rect 34060 17799 34112 17808
rect 34060 17765 34069 17799
rect 34069 17765 34103 17799
rect 34103 17765 34112 17799
rect 34060 17756 34112 17765
rect 31300 17688 31352 17740
rect 32036 17663 32088 17672
rect 32036 17629 32045 17663
rect 32045 17629 32079 17663
rect 32079 17629 32088 17663
rect 32036 17620 32088 17629
rect 33416 17620 33468 17672
rect 33968 17620 34020 17672
rect 18604 17527 18656 17536
rect 18604 17493 18613 17527
rect 18613 17493 18647 17527
rect 18647 17493 18656 17527
rect 18604 17484 18656 17493
rect 18880 17527 18932 17536
rect 18880 17493 18889 17527
rect 18889 17493 18923 17527
rect 18923 17493 18932 17527
rect 18880 17484 18932 17493
rect 18972 17484 19024 17536
rect 29184 17484 29236 17536
rect 30196 17527 30248 17536
rect 30196 17493 30205 17527
rect 30205 17493 30239 17527
rect 30239 17493 30248 17527
rect 30196 17484 30248 17493
rect 31852 17484 31904 17536
rect 33784 17484 33836 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 3424 17323 3476 17332
rect 3424 17289 3433 17323
rect 3433 17289 3467 17323
rect 3467 17289 3476 17323
rect 3424 17280 3476 17289
rect 4252 17323 4304 17332
rect 4252 17289 4261 17323
rect 4261 17289 4295 17323
rect 4295 17289 4304 17323
rect 4252 17280 4304 17289
rect 4068 17212 4120 17264
rect 3240 17187 3292 17196
rect 3240 17153 3249 17187
rect 3249 17153 3283 17187
rect 3283 17153 3292 17187
rect 3240 17144 3292 17153
rect 3792 17076 3844 17128
rect 5724 17280 5776 17332
rect 6368 17280 6420 17332
rect 4804 17212 4856 17264
rect 7748 17280 7800 17332
rect 8484 17144 8536 17196
rect 9496 17280 9548 17332
rect 10140 17280 10192 17332
rect 9404 17212 9456 17264
rect 9680 17212 9732 17264
rect 11152 17280 11204 17332
rect 11980 17323 12032 17332
rect 11980 17289 11989 17323
rect 11989 17289 12023 17323
rect 12023 17289 12032 17323
rect 11980 17280 12032 17289
rect 10324 17212 10376 17264
rect 12256 17280 12308 17332
rect 12440 17280 12492 17332
rect 14004 17323 14056 17332
rect 14004 17289 14013 17323
rect 14013 17289 14047 17323
rect 14047 17289 14056 17323
rect 14004 17280 14056 17289
rect 15568 17280 15620 17332
rect 16212 17280 16264 17332
rect 16764 17280 16816 17332
rect 10416 17187 10468 17196
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 10600 17187 10652 17196
rect 10600 17153 10609 17187
rect 10609 17153 10643 17187
rect 10643 17153 10652 17187
rect 10600 17144 10652 17153
rect 11612 17144 11664 17196
rect 11796 17144 11848 17196
rect 12256 17187 12308 17196
rect 12256 17153 12265 17187
rect 12265 17153 12299 17187
rect 12299 17153 12308 17187
rect 12256 17144 12308 17153
rect 12624 17144 12676 17196
rect 4988 17119 5040 17128
rect 4988 17085 4997 17119
rect 4997 17085 5031 17119
rect 5031 17085 5040 17119
rect 4988 17076 5040 17085
rect 3056 17008 3108 17060
rect 7196 17076 7248 17128
rect 12348 17119 12400 17128
rect 12348 17085 12357 17119
rect 12357 17085 12391 17119
rect 12391 17085 12400 17119
rect 12348 17076 12400 17085
rect 7564 17008 7616 17060
rect 17224 17212 17276 17264
rect 19064 17280 19116 17332
rect 19432 17280 19484 17332
rect 19708 17280 19760 17332
rect 21088 17280 21140 17332
rect 19984 17255 20036 17264
rect 19984 17221 19993 17255
rect 19993 17221 20027 17255
rect 20027 17221 20036 17255
rect 19984 17212 20036 17221
rect 15568 17144 15620 17196
rect 17868 17144 17920 17196
rect 18328 17144 18380 17196
rect 18972 17144 19024 17196
rect 19616 17187 19668 17196
rect 19616 17153 19625 17187
rect 19625 17153 19659 17187
rect 19659 17153 19668 17187
rect 19616 17144 19668 17153
rect 19708 17187 19760 17196
rect 19708 17153 19718 17187
rect 19718 17153 19752 17187
rect 19752 17153 19760 17187
rect 20168 17212 20220 17264
rect 20352 17255 20404 17264
rect 20352 17221 20361 17255
rect 20361 17221 20395 17255
rect 20395 17221 20404 17255
rect 20352 17212 20404 17221
rect 19708 17144 19760 17153
rect 14556 17076 14608 17128
rect 15752 17076 15804 17128
rect 16948 17076 17000 17128
rect 14372 17008 14424 17060
rect 6092 16983 6144 16992
rect 6092 16949 6101 16983
rect 6101 16949 6135 16983
rect 6135 16949 6144 16983
rect 6092 16940 6144 16949
rect 9588 16940 9640 16992
rect 11796 16940 11848 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 18236 16940 18288 16992
rect 18696 16940 18748 16992
rect 20168 17076 20220 17128
rect 20536 17076 20588 17128
rect 20812 17187 20864 17196
rect 23296 17280 23348 17332
rect 23480 17280 23532 17332
rect 28356 17323 28408 17332
rect 28356 17289 28365 17323
rect 28365 17289 28399 17323
rect 28399 17289 28408 17323
rect 28356 17280 28408 17289
rect 20812 17153 20826 17187
rect 20826 17153 20860 17187
rect 20860 17153 20864 17187
rect 20812 17144 20864 17153
rect 19800 16940 19852 16992
rect 20720 17008 20772 17060
rect 22928 17187 22980 17196
rect 22928 17153 22937 17187
rect 22937 17153 22971 17187
rect 22971 17153 22980 17187
rect 22928 17144 22980 17153
rect 27804 17144 27856 17196
rect 29184 17323 29236 17332
rect 29184 17289 29193 17323
rect 29193 17289 29227 17323
rect 29227 17289 29236 17323
rect 29184 17280 29236 17289
rect 30196 17280 30248 17332
rect 28632 17212 28684 17264
rect 32036 17280 32088 17332
rect 32864 17280 32916 17332
rect 33048 17280 33100 17332
rect 33968 17323 34020 17332
rect 33968 17289 33993 17323
rect 33993 17289 34020 17323
rect 33968 17280 34020 17289
rect 23112 17076 23164 17128
rect 29184 17187 29236 17196
rect 29184 17153 29193 17187
rect 29193 17153 29227 17187
rect 29227 17153 29236 17187
rect 29184 17144 29236 17153
rect 29644 17144 29696 17196
rect 31852 17187 31904 17196
rect 31852 17153 31861 17187
rect 31861 17153 31895 17187
rect 31895 17153 31904 17187
rect 31852 17144 31904 17153
rect 32128 17144 32180 17196
rect 33784 17255 33836 17264
rect 33784 17221 33793 17255
rect 33793 17221 33827 17255
rect 33827 17221 33836 17255
rect 33784 17212 33836 17221
rect 32864 17187 32916 17196
rect 32864 17153 32873 17187
rect 32873 17153 32907 17187
rect 32907 17153 32916 17187
rect 32864 17144 32916 17153
rect 34520 17212 34572 17264
rect 23296 17008 23348 17060
rect 25136 17008 25188 17060
rect 28172 17008 28224 17060
rect 24584 16940 24636 16992
rect 28080 16940 28132 16992
rect 30104 17076 30156 17128
rect 32312 17119 32364 17128
rect 32312 17085 32321 17119
rect 32321 17085 32355 17119
rect 32355 17085 32364 17119
rect 32312 17076 32364 17085
rect 32036 17008 32088 17060
rect 29276 16940 29328 16992
rect 29368 16940 29420 16992
rect 30288 16940 30340 16992
rect 31760 16940 31812 16992
rect 31852 16940 31904 16992
rect 32588 17119 32640 17128
rect 32588 17085 32597 17119
rect 32597 17085 32631 17119
rect 32631 17085 32640 17119
rect 32588 17076 32640 17085
rect 34060 17076 34112 17128
rect 34520 17119 34572 17128
rect 34520 17085 34529 17119
rect 34529 17085 34563 17119
rect 34563 17085 34572 17119
rect 34520 17076 34572 17085
rect 33416 16940 33468 16992
rect 34796 16983 34848 16992
rect 34796 16949 34805 16983
rect 34805 16949 34839 16983
rect 34839 16949 34848 16983
rect 34796 16940 34848 16949
rect 35348 16940 35400 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3608 16736 3660 16788
rect 3056 16600 3108 16652
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 2136 16532 2188 16584
rect 1768 16439 1820 16448
rect 1768 16405 1777 16439
rect 1777 16405 1811 16439
rect 1811 16405 1820 16439
rect 1768 16396 1820 16405
rect 1952 16396 2004 16448
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 3148 16396 3200 16448
rect 4252 16464 4304 16516
rect 6092 16736 6144 16788
rect 8484 16668 8536 16720
rect 8300 16600 8352 16652
rect 8852 16600 8904 16652
rect 11980 16668 12032 16720
rect 12256 16668 12308 16720
rect 14280 16736 14332 16788
rect 16580 16736 16632 16788
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 9404 16600 9456 16652
rect 15660 16600 15712 16652
rect 8944 16532 8996 16584
rect 14556 16532 14608 16584
rect 15384 16575 15436 16584
rect 15384 16541 15393 16575
rect 15393 16541 15427 16575
rect 15427 16541 15436 16575
rect 15384 16532 15436 16541
rect 15844 16532 15896 16584
rect 16856 16532 16908 16584
rect 17500 16668 17552 16720
rect 17316 16600 17368 16652
rect 17592 16575 17644 16584
rect 17592 16541 17601 16575
rect 17601 16541 17635 16575
rect 17635 16541 17644 16575
rect 17592 16532 17644 16541
rect 5908 16464 5960 16516
rect 9404 16507 9456 16516
rect 9404 16473 9413 16507
rect 9413 16473 9447 16507
rect 9447 16473 9456 16507
rect 9404 16464 9456 16473
rect 9680 16464 9732 16516
rect 8208 16396 8260 16448
rect 11704 16464 11756 16516
rect 11060 16396 11112 16448
rect 12256 16396 12308 16448
rect 13820 16396 13872 16448
rect 15568 16396 15620 16448
rect 17960 16575 18012 16584
rect 17960 16541 17969 16575
rect 17969 16541 18003 16575
rect 18003 16541 18012 16575
rect 17960 16532 18012 16541
rect 19340 16736 19392 16788
rect 18420 16600 18472 16652
rect 18604 16575 18656 16584
rect 18604 16541 18613 16575
rect 18613 16541 18647 16575
rect 18647 16541 18656 16575
rect 18604 16532 18656 16541
rect 20996 16736 21048 16788
rect 29184 16736 29236 16788
rect 31208 16779 31260 16788
rect 31208 16745 31217 16779
rect 31217 16745 31251 16779
rect 31251 16745 31260 16779
rect 31208 16736 31260 16745
rect 32128 16779 32180 16788
rect 32128 16745 32137 16779
rect 32137 16745 32171 16779
rect 32171 16745 32180 16779
rect 32128 16736 32180 16745
rect 32588 16736 32640 16788
rect 35256 16736 35308 16788
rect 35440 16779 35492 16788
rect 35440 16745 35449 16779
rect 35449 16745 35483 16779
rect 35483 16745 35492 16779
rect 35440 16736 35492 16745
rect 20444 16668 20496 16720
rect 20720 16668 20772 16720
rect 20352 16575 20404 16584
rect 20352 16541 20362 16575
rect 20362 16541 20396 16575
rect 20396 16541 20404 16575
rect 20352 16532 20404 16541
rect 20812 16532 20864 16584
rect 20996 16575 21048 16584
rect 20996 16541 21005 16575
rect 21005 16541 21039 16575
rect 21039 16541 21048 16575
rect 20996 16532 21048 16541
rect 23204 16643 23256 16652
rect 23204 16609 23213 16643
rect 23213 16609 23247 16643
rect 23247 16609 23256 16643
rect 23204 16600 23256 16609
rect 25412 16668 25464 16720
rect 29368 16668 29420 16720
rect 19064 16507 19116 16516
rect 19064 16473 19073 16507
rect 19073 16473 19107 16507
rect 19107 16473 19116 16507
rect 19064 16464 19116 16473
rect 22284 16575 22336 16584
rect 22284 16541 22293 16575
rect 22293 16541 22327 16575
rect 22327 16541 22336 16575
rect 22284 16532 22336 16541
rect 22928 16532 22980 16584
rect 24860 16600 24912 16652
rect 23388 16532 23440 16584
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 26240 16600 26292 16652
rect 26056 16575 26108 16584
rect 16304 16396 16356 16448
rect 16396 16396 16448 16448
rect 16948 16396 17000 16448
rect 18144 16396 18196 16448
rect 18512 16396 18564 16448
rect 22376 16464 22428 16516
rect 22836 16507 22888 16516
rect 22836 16473 22845 16507
rect 22845 16473 22879 16507
rect 22879 16473 22888 16507
rect 22836 16464 22888 16473
rect 23204 16464 23256 16516
rect 23296 16507 23348 16516
rect 23296 16473 23305 16507
rect 23305 16473 23339 16507
rect 23339 16473 23348 16507
rect 23296 16464 23348 16473
rect 20904 16439 20956 16448
rect 20904 16405 20913 16439
rect 20913 16405 20947 16439
rect 20947 16405 20956 16439
rect 20904 16396 20956 16405
rect 23756 16507 23808 16516
rect 23756 16473 23765 16507
rect 23765 16473 23799 16507
rect 23799 16473 23808 16507
rect 23756 16464 23808 16473
rect 26056 16541 26065 16575
rect 26065 16541 26099 16575
rect 26099 16541 26108 16575
rect 26056 16532 26108 16541
rect 32588 16600 32640 16652
rect 35532 16643 35584 16652
rect 35532 16609 35541 16643
rect 35541 16609 35575 16643
rect 35575 16609 35584 16643
rect 35532 16600 35584 16609
rect 30196 16575 30248 16584
rect 30196 16541 30205 16575
rect 30205 16541 30239 16575
rect 30239 16541 30248 16575
rect 30196 16532 30248 16541
rect 30288 16532 30340 16584
rect 30656 16532 30708 16584
rect 30932 16532 30984 16584
rect 31484 16532 31536 16584
rect 31760 16532 31812 16584
rect 25504 16464 25556 16516
rect 29276 16464 29328 16516
rect 25136 16396 25188 16448
rect 26424 16439 26476 16448
rect 26424 16405 26433 16439
rect 26433 16405 26467 16439
rect 26467 16405 26476 16439
rect 26424 16396 26476 16405
rect 28080 16396 28132 16448
rect 30656 16396 30708 16448
rect 30748 16439 30800 16448
rect 30748 16405 30757 16439
rect 30757 16405 30791 16439
rect 30791 16405 30800 16439
rect 30748 16396 30800 16405
rect 32496 16507 32548 16516
rect 32496 16473 32505 16507
rect 32505 16473 32539 16507
rect 32539 16473 32548 16507
rect 32496 16464 32548 16473
rect 34520 16464 34572 16516
rect 34796 16464 34848 16516
rect 35164 16439 35216 16448
rect 35164 16405 35189 16439
rect 35189 16405 35216 16439
rect 35164 16396 35216 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 1400 16192 1452 16244
rect 2964 16192 3016 16244
rect 3608 16192 3660 16244
rect 4620 16192 4672 16244
rect 4988 16192 5040 16244
rect 1952 16124 2004 16176
rect 4804 16124 4856 16176
rect 5448 16192 5500 16244
rect 9404 16192 9456 16244
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 2136 15988 2188 16040
rect 5632 16031 5684 16040
rect 5632 15997 5641 16031
rect 5641 15997 5675 16031
rect 5675 15997 5684 16031
rect 5632 15988 5684 15997
rect 5908 15988 5960 16040
rect 12532 16192 12584 16244
rect 13176 16192 13228 16244
rect 14464 16235 14516 16244
rect 14464 16201 14473 16235
rect 14473 16201 14507 16235
rect 14507 16201 14516 16235
rect 14464 16192 14516 16201
rect 14556 16192 14608 16244
rect 16396 16192 16448 16244
rect 16856 16235 16908 16244
rect 16856 16201 16865 16235
rect 16865 16201 16899 16235
rect 16899 16201 16908 16235
rect 16856 16192 16908 16201
rect 17316 16192 17368 16244
rect 11060 16124 11112 16176
rect 12992 16124 13044 16176
rect 17224 16124 17276 16176
rect 19064 16192 19116 16244
rect 19432 16192 19484 16244
rect 12256 16099 12308 16108
rect 12256 16065 12265 16099
rect 12265 16065 12299 16099
rect 12299 16065 12308 16099
rect 12256 16056 12308 16065
rect 12348 16099 12400 16108
rect 12348 16065 12357 16099
rect 12357 16065 12391 16099
rect 12391 16065 12400 16099
rect 12348 16056 12400 16065
rect 14188 16056 14240 16108
rect 14556 16056 14608 16108
rect 16396 16056 16448 16108
rect 17040 16099 17092 16108
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 18144 16099 18196 16108
rect 18144 16065 18153 16099
rect 18153 16065 18187 16099
rect 18187 16065 18196 16099
rect 18144 16056 18196 16065
rect 18236 16099 18288 16108
rect 18236 16065 18245 16099
rect 18245 16065 18279 16099
rect 18279 16065 18288 16099
rect 18236 16056 18288 16065
rect 18328 16099 18380 16108
rect 18328 16065 18337 16099
rect 18337 16065 18371 16099
rect 18371 16065 18380 16099
rect 18328 16056 18380 16065
rect 18880 16056 18932 16108
rect 10324 16031 10376 16040
rect 10324 15997 10333 16031
rect 10333 15997 10367 16031
rect 10367 15997 10376 16031
rect 10324 15988 10376 15997
rect 11244 15988 11296 16040
rect 11612 15988 11664 16040
rect 12164 15920 12216 15972
rect 13360 15920 13412 15972
rect 15108 15920 15160 15972
rect 3148 15895 3200 15904
rect 3148 15861 3157 15895
rect 3157 15861 3191 15895
rect 3191 15861 3200 15895
rect 3148 15852 3200 15861
rect 3884 15852 3936 15904
rect 16856 15920 16908 15972
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 17132 15920 17184 15972
rect 18328 15852 18380 15904
rect 18604 15895 18656 15904
rect 18604 15861 18613 15895
rect 18613 15861 18647 15895
rect 18647 15861 18656 15895
rect 18604 15852 18656 15861
rect 18696 15852 18748 15904
rect 20444 16124 20496 16176
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 20812 16192 20864 16244
rect 21272 16192 21324 16244
rect 22284 16192 22336 16244
rect 25228 16192 25280 16244
rect 23020 16167 23072 16176
rect 23020 16133 23029 16167
rect 23029 16133 23063 16167
rect 23063 16133 23072 16167
rect 23020 16124 23072 16133
rect 25136 16124 25188 16176
rect 20904 16056 20956 16108
rect 21456 16056 21508 16108
rect 22008 16056 22060 16108
rect 20536 15988 20588 16040
rect 20628 15988 20680 16040
rect 20812 15988 20864 16040
rect 20996 16031 21048 16040
rect 20996 15997 21005 16031
rect 21005 15997 21039 16031
rect 21039 15997 21048 16031
rect 20996 15988 21048 15997
rect 21364 15988 21416 16040
rect 23204 16099 23256 16108
rect 23204 16065 23213 16099
rect 23213 16065 23247 16099
rect 23247 16065 23256 16099
rect 23204 16056 23256 16065
rect 24676 16099 24728 16108
rect 24676 16065 24685 16099
rect 24685 16065 24719 16099
rect 24719 16065 24728 16099
rect 24676 16056 24728 16065
rect 24860 16056 24912 16108
rect 29184 16192 29236 16244
rect 30196 16192 30248 16244
rect 30748 16192 30800 16244
rect 30932 16192 30984 16244
rect 26424 16056 26476 16108
rect 29092 16099 29144 16108
rect 29092 16065 29101 16099
rect 29101 16065 29135 16099
rect 29135 16065 29144 16099
rect 29092 16056 29144 16065
rect 29644 16124 29696 16176
rect 30288 16124 30340 16176
rect 34796 16192 34848 16244
rect 35256 16192 35308 16244
rect 29460 15988 29512 16040
rect 27160 15963 27212 15972
rect 27160 15929 27169 15963
rect 27169 15929 27203 15963
rect 27203 15929 27212 15963
rect 27160 15920 27212 15929
rect 27344 15920 27396 15972
rect 35164 16099 35216 16108
rect 35164 16065 35173 16099
rect 35173 16065 35207 16099
rect 35207 16065 35216 16099
rect 35164 16056 35216 16065
rect 32220 15988 32272 16040
rect 34796 15988 34848 16040
rect 20444 15852 20496 15904
rect 20720 15852 20772 15904
rect 24952 15852 25004 15904
rect 25044 15852 25096 15904
rect 27436 15852 27488 15904
rect 29368 15852 29420 15904
rect 30104 15852 30156 15904
rect 30380 15852 30432 15904
rect 31392 15895 31444 15904
rect 31392 15861 31401 15895
rect 31401 15861 31435 15895
rect 31435 15861 31444 15895
rect 31392 15852 31444 15861
rect 34520 15852 34572 15904
rect 35256 15852 35308 15904
rect 37832 15895 37884 15904
rect 37832 15861 37841 15895
rect 37841 15861 37875 15895
rect 37875 15861 37884 15895
rect 37832 15852 37884 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 940 15648 992 15700
rect 3976 15648 4028 15700
rect 4712 15648 4764 15700
rect 5632 15648 5684 15700
rect 4620 15580 4672 15632
rect 7564 15648 7616 15700
rect 10232 15691 10284 15700
rect 10232 15657 10241 15691
rect 10241 15657 10275 15691
rect 10275 15657 10284 15691
rect 10232 15648 10284 15657
rect 11060 15648 11112 15700
rect 14188 15648 14240 15700
rect 14924 15648 14976 15700
rect 15568 15648 15620 15700
rect 15844 15648 15896 15700
rect 16764 15648 16816 15700
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 3884 15444 3936 15496
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 4160 15487 4212 15496
rect 4160 15453 4169 15487
rect 4169 15453 4203 15487
rect 4203 15453 4212 15487
rect 4160 15444 4212 15453
rect 6184 15555 6236 15564
rect 6184 15521 6193 15555
rect 6193 15521 6227 15555
rect 6227 15521 6236 15555
rect 6184 15512 6236 15521
rect 11244 15512 11296 15564
rect 11612 15580 11664 15632
rect 4804 15444 4856 15496
rect 7840 15444 7892 15496
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 15752 15555 15804 15564
rect 15752 15521 15761 15555
rect 15761 15521 15795 15555
rect 15795 15521 15804 15555
rect 15752 15512 15804 15521
rect 23204 15648 23256 15700
rect 24492 15648 24544 15700
rect 14372 15444 14424 15496
rect 14648 15444 14700 15496
rect 6368 15376 6420 15428
rect 6460 15419 6512 15428
rect 6460 15385 6469 15419
rect 6469 15385 6503 15419
rect 6503 15385 6512 15419
rect 6460 15376 6512 15385
rect 6920 15376 6972 15428
rect 5448 15308 5500 15360
rect 12440 15376 12492 15428
rect 11520 15308 11572 15360
rect 11704 15308 11756 15360
rect 12256 15308 12308 15360
rect 15936 15487 15988 15496
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 17684 15580 17736 15632
rect 18880 15580 18932 15632
rect 18972 15580 19024 15632
rect 16396 15512 16448 15564
rect 16764 15512 16816 15564
rect 16948 15512 17000 15564
rect 17960 15512 18012 15564
rect 18604 15512 18656 15564
rect 15936 15444 15988 15453
rect 15752 15376 15804 15428
rect 18236 15419 18288 15428
rect 18236 15385 18245 15419
rect 18245 15385 18279 15419
rect 18279 15385 18288 15419
rect 18236 15376 18288 15385
rect 18788 15376 18840 15428
rect 19432 15444 19484 15496
rect 21088 15512 21140 15564
rect 22652 15512 22704 15564
rect 20076 15376 20128 15428
rect 18972 15308 19024 15360
rect 19340 15351 19392 15360
rect 19340 15317 19349 15351
rect 19349 15317 19383 15351
rect 19383 15317 19392 15351
rect 19340 15308 19392 15317
rect 19984 15308 20036 15360
rect 20536 15308 20588 15360
rect 22008 15444 22060 15496
rect 23020 15444 23072 15496
rect 23940 15444 23992 15496
rect 24492 15487 24544 15496
rect 24492 15453 24501 15487
rect 24501 15453 24535 15487
rect 24535 15453 24544 15487
rect 24492 15444 24544 15453
rect 24676 15444 24728 15496
rect 25228 15487 25280 15496
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 27344 15648 27396 15700
rect 29460 15648 29512 15700
rect 30748 15648 30800 15700
rect 31392 15648 31444 15700
rect 32220 15648 32272 15700
rect 32588 15648 32640 15700
rect 32864 15648 32916 15700
rect 34796 15648 34848 15700
rect 35532 15648 35584 15700
rect 27160 15512 27212 15564
rect 27436 15512 27488 15564
rect 25504 15444 25556 15496
rect 26056 15444 26108 15496
rect 26240 15444 26292 15496
rect 27068 15444 27120 15496
rect 27436 15376 27488 15428
rect 24676 15308 24728 15360
rect 25504 15308 25556 15360
rect 25688 15308 25740 15360
rect 27344 15308 27396 15360
rect 28080 15444 28132 15496
rect 29092 15444 29144 15496
rect 34796 15555 34848 15564
rect 34796 15521 34805 15555
rect 34805 15521 34839 15555
rect 34839 15521 34848 15555
rect 34796 15512 34848 15521
rect 35624 15555 35676 15564
rect 35624 15521 35633 15555
rect 35633 15521 35667 15555
rect 35667 15521 35676 15555
rect 35624 15512 35676 15521
rect 32864 15444 32916 15496
rect 33416 15487 33468 15496
rect 33416 15453 33425 15487
rect 33425 15453 33459 15487
rect 33459 15453 33468 15487
rect 33416 15444 33468 15453
rect 34612 15444 34664 15496
rect 34704 15444 34756 15496
rect 30288 15376 30340 15428
rect 32220 15376 32272 15428
rect 28356 15351 28408 15360
rect 28356 15317 28365 15351
rect 28365 15317 28399 15351
rect 28399 15317 28408 15351
rect 28356 15308 28408 15317
rect 30656 15351 30708 15360
rect 30656 15317 30665 15351
rect 30665 15317 30699 15351
rect 30699 15317 30708 15351
rect 30656 15308 30708 15317
rect 32588 15351 32640 15360
rect 32588 15317 32597 15351
rect 32597 15317 32631 15351
rect 32631 15317 32640 15351
rect 32588 15308 32640 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 5448 15104 5500 15156
rect 6460 15104 6512 15156
rect 7564 15147 7616 15156
rect 7564 15113 7573 15147
rect 7573 15113 7607 15147
rect 7607 15113 7616 15147
rect 7564 15104 7616 15113
rect 8300 15104 8352 15156
rect 8760 15104 8812 15156
rect 9496 15104 9548 15156
rect 12164 15104 12216 15156
rect 12440 15104 12492 15156
rect 14556 15104 14608 15156
rect 14924 15104 14976 15156
rect 16396 15104 16448 15156
rect 18788 15104 18840 15156
rect 26056 15104 26108 15156
rect 27344 15104 27396 15156
rect 27620 15104 27672 15156
rect 27896 15104 27948 15156
rect 32588 15104 32640 15156
rect 34796 15104 34848 15156
rect 3240 14968 3292 15020
rect 4160 15036 4212 15088
rect 3976 14968 4028 15020
rect 3148 14943 3200 14952
rect 3148 14909 3157 14943
rect 3157 14909 3191 14943
rect 3191 14909 3200 14943
rect 3148 14900 3200 14909
rect 4252 14943 4304 14952
rect 4252 14909 4261 14943
rect 4261 14909 4295 14943
rect 4295 14909 4304 14943
rect 4252 14900 4304 14909
rect 4068 14832 4120 14884
rect 2504 14807 2556 14816
rect 2504 14773 2513 14807
rect 2513 14773 2547 14807
rect 2547 14773 2556 14807
rect 2504 14764 2556 14773
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 3884 14764 3936 14816
rect 4620 15036 4672 15088
rect 4712 15011 4764 15020
rect 4712 14977 4721 15011
rect 4721 14977 4755 15011
rect 4755 14977 4764 15011
rect 4712 14968 4764 14977
rect 7196 14900 7248 14952
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 8944 14968 8996 15020
rect 9588 15036 9640 15088
rect 10784 15036 10836 15088
rect 9496 14943 9548 14952
rect 9496 14909 9505 14943
rect 9505 14909 9539 14943
rect 9539 14909 9548 14943
rect 9496 14900 9548 14909
rect 8116 14832 8168 14884
rect 9036 14875 9088 14884
rect 9036 14841 9045 14875
rect 9045 14841 9079 14875
rect 9079 14841 9088 14875
rect 9036 14832 9088 14841
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 13728 14968 13780 15020
rect 13820 14968 13872 15020
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 14372 14968 14424 15020
rect 12624 14900 12676 14952
rect 12808 14900 12860 14952
rect 14648 14900 14700 14952
rect 14280 14832 14332 14884
rect 15016 14900 15068 14952
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 15936 14968 15988 15020
rect 16120 14968 16172 15020
rect 16212 15011 16264 15020
rect 16212 14977 16221 15011
rect 16221 14977 16255 15011
rect 16255 14977 16264 15011
rect 16212 14968 16264 14977
rect 16948 14968 17000 15020
rect 17040 15011 17092 15020
rect 17040 14977 17049 15011
rect 17049 14977 17083 15011
rect 17083 14977 17092 15011
rect 17040 14968 17092 14977
rect 16304 14900 16356 14952
rect 17224 14968 17276 15020
rect 17684 15011 17736 15020
rect 17684 14977 17693 15011
rect 17693 14977 17727 15011
rect 17727 14977 17736 15011
rect 17684 14968 17736 14977
rect 18604 14968 18656 15020
rect 20444 15036 20496 15088
rect 19432 14968 19484 15020
rect 19984 14968 20036 15020
rect 20168 15011 20220 15020
rect 20168 14977 20177 15011
rect 20177 14977 20211 15011
rect 20211 14977 20220 15011
rect 20168 14968 20220 14977
rect 18236 14900 18288 14952
rect 20812 14968 20864 15020
rect 23204 15011 23256 15020
rect 23204 14977 23213 15011
rect 23213 14977 23247 15011
rect 23247 14977 23256 15011
rect 23204 14968 23256 14977
rect 25688 15011 25740 15020
rect 25688 14977 25697 15011
rect 25697 14977 25731 15011
rect 25731 14977 25740 15011
rect 25688 14968 25740 14977
rect 21824 14943 21876 14952
rect 21824 14909 21833 14943
rect 21833 14909 21867 14943
rect 21867 14909 21876 14943
rect 21824 14900 21876 14909
rect 22100 14900 22152 14952
rect 26332 14968 26384 15020
rect 26424 14968 26476 15020
rect 27160 14968 27212 15020
rect 27804 15011 27856 15020
rect 27804 14977 27813 15011
rect 27813 14977 27847 15011
rect 27847 14977 27856 15011
rect 27804 14968 27856 14977
rect 26148 14900 26200 14952
rect 28172 14900 28224 14952
rect 28448 15011 28500 15020
rect 28448 14977 28457 15011
rect 28457 14977 28491 15011
rect 28491 14977 28500 15011
rect 28448 14968 28500 14977
rect 28724 14968 28776 15020
rect 8668 14807 8720 14816
rect 8668 14773 8677 14807
rect 8677 14773 8711 14807
rect 8711 14773 8720 14807
rect 8668 14764 8720 14773
rect 8944 14764 8996 14816
rect 9772 14807 9824 14816
rect 9772 14773 9781 14807
rect 9781 14773 9815 14807
rect 9815 14773 9824 14807
rect 9772 14764 9824 14773
rect 10232 14764 10284 14816
rect 11980 14764 12032 14816
rect 18788 14875 18840 14884
rect 18788 14841 18797 14875
rect 18797 14841 18831 14875
rect 18831 14841 18840 14875
rect 18788 14832 18840 14841
rect 19432 14832 19484 14884
rect 24124 14832 24176 14884
rect 24768 14832 24820 14884
rect 16396 14807 16448 14816
rect 16396 14773 16405 14807
rect 16405 14773 16439 14807
rect 16439 14773 16448 14807
rect 16396 14764 16448 14773
rect 17684 14764 17736 14816
rect 20536 14807 20588 14816
rect 20536 14773 20545 14807
rect 20545 14773 20579 14807
rect 20579 14773 20588 14807
rect 20536 14764 20588 14773
rect 20812 14764 20864 14816
rect 22192 14764 22244 14816
rect 22284 14764 22336 14816
rect 24584 14764 24636 14816
rect 25596 14807 25648 14816
rect 25596 14773 25605 14807
rect 25605 14773 25639 14807
rect 25639 14773 25648 14807
rect 25596 14764 25648 14773
rect 26332 14764 26384 14816
rect 28448 14832 28500 14884
rect 28540 14832 28592 14884
rect 30656 15011 30708 15020
rect 30656 14977 30665 15011
rect 30665 14977 30699 15011
rect 30699 14977 30708 15011
rect 30656 14968 30708 14977
rect 30840 15011 30892 15020
rect 30840 14977 30849 15011
rect 30849 14977 30883 15011
rect 30883 14977 30892 15011
rect 30840 14968 30892 14977
rect 29920 14900 29972 14952
rect 30564 14900 30616 14952
rect 31116 15011 31168 15020
rect 31116 14977 31125 15011
rect 31125 14977 31159 15011
rect 31159 14977 31168 15011
rect 31116 14968 31168 14977
rect 33048 15011 33100 15020
rect 33048 14977 33057 15011
rect 33057 14977 33091 15011
rect 33091 14977 33100 15011
rect 33048 14968 33100 14977
rect 32956 14943 33008 14952
rect 32956 14909 32965 14943
rect 32965 14909 32999 14943
rect 32999 14909 33008 14943
rect 32956 14900 33008 14909
rect 30472 14832 30524 14884
rect 30748 14832 30800 14884
rect 28816 14764 28868 14816
rect 31024 14807 31076 14816
rect 31024 14773 31033 14807
rect 31033 14773 31067 14807
rect 31067 14773 31076 14807
rect 31024 14764 31076 14773
rect 31392 14764 31444 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3240 14560 3292 14612
rect 3608 14560 3660 14612
rect 4068 14603 4120 14612
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 7472 14560 7524 14612
rect 14096 14560 14148 14612
rect 15844 14560 15896 14612
rect 17040 14603 17092 14612
rect 17040 14569 17049 14603
rect 17049 14569 17083 14603
rect 17083 14569 17092 14603
rect 17040 14560 17092 14569
rect 17408 14603 17460 14612
rect 17408 14569 17417 14603
rect 17417 14569 17451 14603
rect 17451 14569 17460 14603
rect 17408 14560 17460 14569
rect 22284 14603 22336 14612
rect 22284 14569 22293 14603
rect 22293 14569 22327 14603
rect 22327 14569 22336 14603
rect 22284 14560 22336 14569
rect 23112 14560 23164 14612
rect 26424 14560 26476 14612
rect 28356 14560 28408 14612
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 13820 14492 13872 14544
rect 3700 14424 3752 14476
rect 4620 14356 4672 14408
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 8576 14424 8628 14476
rect 9036 14356 9088 14408
rect 9220 14399 9272 14408
rect 9220 14365 9229 14399
rect 9229 14365 9263 14399
rect 9263 14365 9272 14399
rect 9220 14356 9272 14365
rect 10232 14424 10284 14476
rect 12164 14424 12216 14476
rect 12624 14424 12676 14476
rect 14372 14424 14424 14476
rect 15016 14424 15068 14476
rect 17776 14492 17828 14544
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 1676 14331 1728 14340
rect 1676 14297 1685 14331
rect 1685 14297 1719 14331
rect 1719 14297 1728 14331
rect 1676 14288 1728 14297
rect 2964 14288 3016 14340
rect 5908 14331 5960 14340
rect 5908 14297 5917 14331
rect 5917 14297 5951 14331
rect 5951 14297 5960 14331
rect 5908 14288 5960 14297
rect 6920 14288 6972 14340
rect 9588 14331 9640 14340
rect 9588 14297 9597 14331
rect 9597 14297 9631 14331
rect 9631 14297 9640 14331
rect 9588 14288 9640 14297
rect 12256 14288 12308 14340
rect 8668 14220 8720 14272
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 16396 14356 16448 14408
rect 16672 14356 16724 14408
rect 16764 14399 16816 14408
rect 16764 14365 16773 14399
rect 16773 14365 16807 14399
rect 16807 14365 16816 14399
rect 16764 14356 16816 14365
rect 16948 14288 17000 14340
rect 14004 14220 14056 14272
rect 14280 14220 14332 14272
rect 15752 14220 15804 14272
rect 15936 14220 15988 14272
rect 17684 14424 17736 14476
rect 17408 14288 17460 14340
rect 20168 14492 20220 14544
rect 20536 14492 20588 14544
rect 20628 14492 20680 14544
rect 20076 14356 20128 14408
rect 20444 14288 20496 14340
rect 21088 14356 21140 14408
rect 22744 14492 22796 14544
rect 29184 14492 29236 14544
rect 31024 14492 31076 14544
rect 22100 14424 22152 14476
rect 22284 14424 22336 14476
rect 23204 14424 23256 14476
rect 21824 14288 21876 14340
rect 22836 14356 22888 14408
rect 30656 14424 30708 14476
rect 30840 14424 30892 14476
rect 23480 14356 23532 14408
rect 23204 14288 23256 14340
rect 24124 14356 24176 14408
rect 25504 14356 25556 14408
rect 27160 14356 27212 14408
rect 31576 14492 31628 14544
rect 31668 14424 31720 14476
rect 32956 14560 33008 14612
rect 30748 14288 30800 14340
rect 19340 14220 19392 14272
rect 19984 14220 20036 14272
rect 22836 14220 22888 14272
rect 25136 14220 25188 14272
rect 25780 14220 25832 14272
rect 26240 14220 26292 14272
rect 27068 14220 27120 14272
rect 29276 14220 29328 14272
rect 30196 14220 30248 14272
rect 30380 14220 30432 14272
rect 31208 14220 31260 14272
rect 31392 14220 31444 14272
rect 33784 14220 33836 14272
rect 34060 14220 34112 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1676 14016 1728 14068
rect 2504 14016 2556 14068
rect 5908 14016 5960 14068
rect 8668 14059 8720 14068
rect 8668 14025 8677 14059
rect 8677 14025 8711 14059
rect 8711 14025 8720 14059
rect 8668 14016 8720 14025
rect 11980 14016 12032 14068
rect 13820 14016 13872 14068
rect 16948 14016 17000 14068
rect 19432 14016 19484 14068
rect 21088 14016 21140 14068
rect 21272 14016 21324 14068
rect 22192 14016 22244 14068
rect 22836 14059 22888 14068
rect 22836 14025 22845 14059
rect 22845 14025 22879 14059
rect 22879 14025 22888 14059
rect 22836 14016 22888 14025
rect 7472 13948 7524 14000
rect 8300 13948 8352 14000
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 10140 13948 10192 14000
rect 9956 13880 10008 13932
rect 12808 13880 12860 13932
rect 13360 13880 13412 13932
rect 14648 13923 14700 13932
rect 14648 13889 14657 13923
rect 14657 13889 14691 13923
rect 14691 13889 14700 13923
rect 14648 13880 14700 13889
rect 15200 13880 15252 13932
rect 17316 13948 17368 14000
rect 20076 13948 20128 14000
rect 17132 13880 17184 13932
rect 17408 13880 17460 13932
rect 5540 13812 5592 13864
rect 7196 13855 7248 13864
rect 7196 13821 7205 13855
rect 7205 13821 7239 13855
rect 7239 13821 7248 13855
rect 7196 13812 7248 13821
rect 16856 13812 16908 13864
rect 19616 13880 19668 13932
rect 19708 13923 19760 13932
rect 19708 13889 19717 13923
rect 19717 13889 19751 13923
rect 19751 13889 19760 13923
rect 19708 13880 19760 13889
rect 10968 13744 11020 13796
rect 18420 13744 18472 13796
rect 19156 13744 19208 13796
rect 9404 13676 9456 13728
rect 12532 13676 12584 13728
rect 15568 13676 15620 13728
rect 17408 13719 17460 13728
rect 17408 13685 17417 13719
rect 17417 13685 17451 13719
rect 17451 13685 17460 13719
rect 17408 13676 17460 13685
rect 17868 13676 17920 13728
rect 19432 13676 19484 13728
rect 20536 13948 20588 14000
rect 20444 13880 20496 13932
rect 20720 13880 20772 13932
rect 23204 13948 23256 14000
rect 21824 13880 21876 13932
rect 24124 13923 24176 13932
rect 24124 13889 24133 13923
rect 24133 13889 24167 13923
rect 24167 13889 24176 13923
rect 24124 13880 24176 13889
rect 24768 13923 24820 13932
rect 24768 13889 24777 13923
rect 24777 13889 24811 13923
rect 24811 13889 24820 13923
rect 24768 13880 24820 13889
rect 25044 13923 25096 13932
rect 25044 13889 25053 13923
rect 25053 13889 25087 13923
rect 25087 13889 25096 13923
rect 25044 13880 25096 13889
rect 25136 13923 25188 13932
rect 25136 13889 25145 13923
rect 25145 13889 25179 13923
rect 25179 13889 25188 13923
rect 25136 13880 25188 13889
rect 25780 13948 25832 14000
rect 26332 14016 26384 14068
rect 21364 13744 21416 13796
rect 22376 13812 22428 13864
rect 22560 13812 22612 13864
rect 22744 13812 22796 13864
rect 22928 13744 22980 13796
rect 23204 13855 23256 13864
rect 23204 13821 23213 13855
rect 23213 13821 23247 13855
rect 23247 13821 23256 13855
rect 23204 13812 23256 13821
rect 22560 13676 22612 13728
rect 22744 13676 22796 13728
rect 23480 13812 23532 13864
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 23848 13812 23900 13864
rect 26148 13880 26200 13932
rect 27252 14016 27304 14068
rect 28448 14016 28500 14068
rect 29184 14016 29236 14068
rect 30840 14016 30892 14068
rect 31484 14016 31536 14068
rect 32864 14059 32916 14068
rect 32864 14025 32873 14059
rect 32873 14025 32907 14059
rect 32907 14025 32916 14059
rect 32864 14016 32916 14025
rect 27068 13923 27120 13932
rect 27068 13889 27077 13923
rect 27077 13889 27111 13923
rect 27111 13889 27120 13923
rect 27068 13880 27120 13889
rect 27804 13948 27856 14000
rect 28080 13880 28132 13932
rect 28816 13923 28868 13932
rect 28816 13889 28825 13923
rect 28825 13889 28859 13923
rect 28859 13889 28868 13923
rect 28816 13880 28868 13889
rect 24400 13787 24452 13796
rect 24400 13753 24409 13787
rect 24409 13753 24443 13787
rect 24443 13753 24452 13787
rect 24400 13744 24452 13753
rect 25504 13744 25556 13796
rect 24216 13676 24268 13728
rect 29000 13812 29052 13864
rect 27252 13744 27304 13796
rect 29184 13880 29236 13932
rect 30104 13812 30156 13864
rect 30380 13923 30432 13932
rect 30380 13889 30389 13923
rect 30389 13889 30423 13923
rect 30423 13889 30432 13923
rect 30380 13880 30432 13889
rect 30840 13880 30892 13932
rect 30472 13855 30524 13864
rect 30472 13821 30481 13855
rect 30481 13821 30515 13855
rect 30515 13821 30524 13855
rect 30472 13812 30524 13821
rect 25780 13676 25832 13728
rect 26240 13676 26292 13728
rect 26700 13676 26752 13728
rect 27160 13719 27212 13728
rect 27160 13685 27169 13719
rect 27169 13685 27203 13719
rect 27203 13685 27212 13719
rect 27160 13676 27212 13685
rect 28540 13719 28592 13728
rect 28540 13685 28549 13719
rect 28549 13685 28583 13719
rect 28583 13685 28592 13719
rect 28540 13676 28592 13685
rect 29276 13744 29328 13796
rect 30748 13744 30800 13796
rect 32404 13812 32456 13864
rect 32956 13923 33008 13932
rect 32956 13889 32965 13923
rect 32965 13889 32999 13923
rect 32999 13889 33008 13923
rect 32956 13880 33008 13889
rect 33232 13923 33284 13932
rect 33232 13889 33241 13923
rect 33241 13889 33275 13923
rect 33275 13889 33284 13923
rect 33232 13880 33284 13889
rect 33508 13880 33560 13932
rect 29460 13676 29512 13728
rect 31852 13719 31904 13728
rect 31852 13685 31861 13719
rect 31861 13685 31895 13719
rect 31895 13685 31904 13719
rect 31852 13676 31904 13685
rect 32588 13676 32640 13728
rect 33140 13676 33192 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 9036 13472 9088 13524
rect 10324 13472 10376 13524
rect 10416 13472 10468 13524
rect 1400 13336 1452 13388
rect 5632 13336 5684 13388
rect 6276 13336 6328 13388
rect 3332 13268 3384 13320
rect 3792 13268 3844 13320
rect 3976 13200 4028 13252
rect 4620 13243 4672 13252
rect 4620 13209 4629 13243
rect 4629 13209 4663 13243
rect 4663 13209 4672 13243
rect 4620 13200 4672 13209
rect 2964 13132 3016 13184
rect 6920 13336 6972 13388
rect 7196 13379 7248 13388
rect 7196 13345 7205 13379
rect 7205 13345 7239 13379
rect 7239 13345 7248 13379
rect 7196 13336 7248 13345
rect 9588 13336 9640 13388
rect 9220 13268 9272 13320
rect 9956 13243 10008 13252
rect 9956 13209 9965 13243
rect 9965 13209 9999 13243
rect 9999 13209 10008 13243
rect 9956 13200 10008 13209
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 11244 13472 11296 13524
rect 11888 13336 11940 13388
rect 13820 13472 13872 13524
rect 14740 13472 14792 13524
rect 15292 13472 15344 13524
rect 16764 13472 16816 13524
rect 17224 13472 17276 13524
rect 17868 13515 17920 13524
rect 17868 13481 17877 13515
rect 17877 13481 17911 13515
rect 17911 13481 17920 13515
rect 17868 13472 17920 13481
rect 18420 13515 18472 13524
rect 18420 13481 18429 13515
rect 18429 13481 18463 13515
rect 18463 13481 18472 13515
rect 18420 13472 18472 13481
rect 12624 13336 12676 13388
rect 13360 13336 13412 13388
rect 16856 13404 16908 13456
rect 12532 13268 12584 13320
rect 11152 13200 11204 13252
rect 6552 13175 6604 13184
rect 6552 13141 6561 13175
rect 6561 13141 6595 13175
rect 6595 13141 6604 13175
rect 6552 13132 6604 13141
rect 8024 13132 8076 13184
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 9496 13175 9548 13184
rect 9496 13141 9505 13175
rect 9505 13141 9539 13175
rect 9539 13141 9548 13175
rect 9496 13132 9548 13141
rect 9588 13175 9640 13184
rect 9588 13141 9597 13175
rect 9597 13141 9631 13175
rect 9631 13141 9640 13175
rect 9588 13132 9640 13141
rect 12256 13200 12308 13252
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 13728 13200 13780 13252
rect 14648 13200 14700 13252
rect 15200 13243 15252 13252
rect 15200 13209 15209 13243
rect 15209 13209 15243 13243
rect 15243 13209 15252 13243
rect 15200 13200 15252 13209
rect 16672 13243 16724 13252
rect 16672 13209 16681 13243
rect 16681 13209 16715 13243
rect 16715 13209 16724 13243
rect 16672 13200 16724 13209
rect 13636 13175 13688 13184
rect 13636 13141 13645 13175
rect 13645 13141 13679 13175
rect 13679 13141 13688 13175
rect 13636 13132 13688 13141
rect 13820 13132 13872 13184
rect 15292 13132 15344 13184
rect 15568 13132 15620 13184
rect 18328 13200 18380 13252
rect 19708 13515 19760 13524
rect 19708 13481 19717 13515
rect 19717 13481 19751 13515
rect 19751 13481 19760 13515
rect 19708 13472 19760 13481
rect 20628 13515 20680 13524
rect 19340 13404 19392 13456
rect 18696 13268 18748 13320
rect 19616 13268 19668 13320
rect 20628 13481 20637 13515
rect 20637 13481 20671 13515
rect 20671 13481 20680 13515
rect 20628 13472 20680 13481
rect 20444 13404 20496 13456
rect 21824 13404 21876 13456
rect 22744 13404 22796 13456
rect 22928 13447 22980 13456
rect 22928 13413 22937 13447
rect 22937 13413 22971 13447
rect 22971 13413 22980 13447
rect 22928 13404 22980 13413
rect 23848 13404 23900 13456
rect 20076 13311 20128 13320
rect 20076 13277 20085 13311
rect 20085 13277 20119 13311
rect 20119 13277 20128 13311
rect 20076 13268 20128 13277
rect 19156 13200 19208 13252
rect 20536 13268 20588 13320
rect 21088 13311 21140 13320
rect 21088 13277 21097 13311
rect 21097 13277 21131 13311
rect 21131 13277 21140 13311
rect 21088 13268 21140 13277
rect 21364 13311 21416 13320
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 22376 13311 22428 13320
rect 22376 13277 22385 13311
rect 22385 13277 22419 13311
rect 22419 13277 22428 13311
rect 22376 13268 22428 13277
rect 23204 13311 23256 13320
rect 23204 13277 23213 13311
rect 23213 13277 23247 13311
rect 23247 13277 23256 13311
rect 23204 13268 23256 13277
rect 24124 13268 24176 13320
rect 25780 13336 25832 13388
rect 26240 13379 26292 13388
rect 24860 13268 24912 13320
rect 25596 13268 25648 13320
rect 25872 13311 25924 13320
rect 25872 13277 25881 13311
rect 25881 13277 25915 13311
rect 25915 13277 25924 13311
rect 25872 13268 25924 13277
rect 18696 13175 18748 13184
rect 18696 13141 18705 13175
rect 18705 13141 18739 13175
rect 18739 13141 18748 13175
rect 18696 13132 18748 13141
rect 20168 13132 20220 13184
rect 20536 13132 20588 13184
rect 24492 13200 24544 13252
rect 25504 13200 25556 13252
rect 26240 13345 26249 13379
rect 26249 13345 26283 13379
rect 26283 13345 26292 13379
rect 26240 13336 26292 13345
rect 26976 13404 27028 13456
rect 27804 13472 27856 13524
rect 28172 13472 28224 13524
rect 29000 13472 29052 13524
rect 29184 13515 29236 13524
rect 29184 13481 29193 13515
rect 29193 13481 29227 13515
rect 29227 13481 29236 13515
rect 29184 13472 29236 13481
rect 32404 13472 32456 13524
rect 33232 13515 33284 13524
rect 33232 13481 33241 13515
rect 33241 13481 33275 13515
rect 33275 13481 33284 13515
rect 33232 13472 33284 13481
rect 33416 13472 33468 13524
rect 28356 13404 28408 13456
rect 30288 13404 30340 13456
rect 31208 13404 31260 13456
rect 32128 13404 32180 13456
rect 26516 13311 26568 13320
rect 26516 13277 26525 13311
rect 26525 13277 26559 13311
rect 26559 13277 26568 13311
rect 26516 13268 26568 13277
rect 26792 13311 26844 13320
rect 26792 13277 26801 13311
rect 26801 13277 26835 13311
rect 26835 13277 26844 13311
rect 26792 13268 26844 13277
rect 27068 13311 27120 13320
rect 27068 13277 27077 13311
rect 27077 13277 27111 13311
rect 27111 13277 27120 13311
rect 27068 13268 27120 13277
rect 27160 13311 27212 13320
rect 27160 13277 27169 13311
rect 27169 13277 27203 13311
rect 27203 13277 27212 13311
rect 27160 13268 27212 13277
rect 21180 13132 21232 13184
rect 21548 13175 21600 13184
rect 21548 13141 21557 13175
rect 21557 13141 21591 13175
rect 21591 13141 21600 13175
rect 21548 13132 21600 13141
rect 22192 13132 22244 13184
rect 26700 13200 26752 13252
rect 25780 13175 25832 13184
rect 25780 13141 25789 13175
rect 25789 13141 25823 13175
rect 25823 13141 25832 13175
rect 25780 13132 25832 13141
rect 26516 13132 26568 13184
rect 28540 13311 28592 13320
rect 28540 13277 28549 13311
rect 28549 13277 28583 13311
rect 28583 13277 28592 13311
rect 28540 13268 28592 13277
rect 29276 13311 29328 13320
rect 29276 13277 29285 13311
rect 29285 13277 29319 13311
rect 29319 13277 29328 13311
rect 29276 13268 29328 13277
rect 29460 13268 29512 13320
rect 31208 13268 31260 13320
rect 32864 13311 32916 13320
rect 32864 13277 32873 13311
rect 32873 13277 32907 13311
rect 32907 13277 32916 13311
rect 32864 13268 32916 13277
rect 33140 13268 33192 13320
rect 31300 13200 31352 13252
rect 31668 13200 31720 13252
rect 32588 13243 32640 13252
rect 32588 13209 32597 13243
rect 32597 13209 32631 13243
rect 32631 13209 32640 13243
rect 32588 13200 32640 13209
rect 33508 13311 33560 13320
rect 33508 13277 33517 13311
rect 33517 13277 33551 13311
rect 33551 13277 33560 13311
rect 33508 13268 33560 13277
rect 33876 13311 33928 13320
rect 33876 13277 33885 13311
rect 33885 13277 33919 13311
rect 33919 13277 33928 13311
rect 33876 13268 33928 13277
rect 28448 13132 28500 13184
rect 28908 13132 28960 13184
rect 29644 13175 29696 13184
rect 29644 13141 29653 13175
rect 29653 13141 29687 13175
rect 29687 13141 29696 13175
rect 29644 13132 29696 13141
rect 32956 13132 33008 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 3976 12928 4028 12980
rect 4620 12928 4672 12980
rect 6552 12928 6604 12980
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 2964 12792 3016 12844
rect 3976 12835 4028 12844
rect 3976 12801 3985 12835
rect 3985 12801 4019 12835
rect 4019 12801 4028 12835
rect 3976 12792 4028 12801
rect 4436 12835 4488 12844
rect 4436 12801 4445 12835
rect 4445 12801 4479 12835
rect 4479 12801 4488 12835
rect 4436 12792 4488 12801
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 3884 12724 3936 12776
rect 3792 12656 3844 12708
rect 4712 12792 4764 12844
rect 5816 12792 5868 12844
rect 6920 12860 6972 12912
rect 6368 12835 6420 12844
rect 6368 12801 6377 12835
rect 6377 12801 6411 12835
rect 6411 12801 6420 12835
rect 6368 12792 6420 12801
rect 8024 12928 8076 12980
rect 9864 12928 9916 12980
rect 10416 12928 10468 12980
rect 13636 12928 13688 12980
rect 13820 12928 13872 12980
rect 15200 12928 15252 12980
rect 20076 12928 20128 12980
rect 21180 12928 21232 12980
rect 21732 12928 21784 12980
rect 8576 12903 8628 12912
rect 8576 12869 8585 12903
rect 8585 12869 8619 12903
rect 8619 12869 8628 12903
rect 8576 12860 8628 12869
rect 9680 12792 9732 12844
rect 10232 12792 10284 12844
rect 19248 12860 19300 12912
rect 9588 12656 9640 12708
rect 11888 12792 11940 12844
rect 11980 12724 12032 12776
rect 12716 12792 12768 12844
rect 14924 12792 14976 12844
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 15476 12792 15528 12801
rect 13176 12767 13228 12776
rect 13176 12733 13185 12767
rect 13185 12733 13219 12767
rect 13219 12733 13228 12767
rect 13176 12724 13228 12733
rect 15660 12767 15712 12776
rect 15660 12733 15669 12767
rect 15669 12733 15703 12767
rect 15703 12733 15712 12767
rect 15660 12724 15712 12733
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 20168 12835 20220 12844
rect 20168 12801 20177 12835
rect 20177 12801 20211 12835
rect 20211 12801 20220 12835
rect 20168 12792 20220 12801
rect 20996 12860 21048 12912
rect 21548 12860 21600 12912
rect 24768 12928 24820 12980
rect 25872 12928 25924 12980
rect 26700 12928 26752 12980
rect 29644 12928 29696 12980
rect 31208 12971 31260 12980
rect 31208 12937 31217 12971
rect 31217 12937 31251 12971
rect 31251 12937 31260 12971
rect 31208 12928 31260 12937
rect 19984 12724 20036 12776
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 21824 12835 21876 12844
rect 21824 12801 21833 12835
rect 21833 12801 21867 12835
rect 21867 12801 21876 12835
rect 21824 12792 21876 12801
rect 3056 12588 3108 12640
rect 10140 12631 10192 12640
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 10140 12588 10192 12597
rect 15108 12631 15160 12640
rect 15108 12597 15117 12631
rect 15117 12597 15151 12631
rect 15151 12597 15160 12631
rect 15108 12588 15160 12597
rect 16396 12588 16448 12640
rect 19432 12588 19484 12640
rect 19892 12631 19944 12640
rect 19892 12597 19901 12631
rect 19901 12597 19935 12631
rect 19935 12597 19944 12631
rect 19892 12588 19944 12597
rect 20628 12588 20680 12640
rect 21364 12588 21416 12640
rect 22192 12767 22244 12776
rect 22192 12733 22201 12767
rect 22201 12733 22235 12767
rect 22235 12733 22244 12767
rect 22192 12724 22244 12733
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 23204 12792 23256 12844
rect 24216 12792 24268 12844
rect 24124 12724 24176 12776
rect 24308 12724 24360 12776
rect 24492 12767 24544 12776
rect 24492 12733 24501 12767
rect 24501 12733 24535 12767
rect 24535 12733 24544 12767
rect 24492 12724 24544 12733
rect 25596 12792 25648 12844
rect 26332 12792 26384 12844
rect 22560 12656 22612 12708
rect 25228 12767 25280 12776
rect 25228 12733 25237 12767
rect 25237 12733 25271 12767
rect 25271 12733 25280 12767
rect 25228 12724 25280 12733
rect 26516 12835 26568 12844
rect 26516 12801 26525 12835
rect 26525 12801 26559 12835
rect 26559 12801 26568 12835
rect 26516 12792 26568 12801
rect 31852 12971 31904 12980
rect 31852 12937 31861 12971
rect 31861 12937 31895 12971
rect 31895 12937 31904 12971
rect 31852 12928 31904 12937
rect 32864 12971 32916 12980
rect 32864 12937 32873 12971
rect 32873 12937 32907 12971
rect 32907 12937 32916 12971
rect 32864 12928 32916 12937
rect 33140 12928 33192 12980
rect 26884 12724 26936 12776
rect 28172 12724 28224 12776
rect 30012 12792 30064 12844
rect 30380 12792 30432 12844
rect 30656 12835 30708 12844
rect 30656 12801 30665 12835
rect 30665 12801 30699 12835
rect 30699 12801 30708 12835
rect 30656 12792 30708 12801
rect 31208 12835 31260 12844
rect 31208 12801 31217 12835
rect 31217 12801 31251 12835
rect 31251 12801 31260 12835
rect 31208 12792 31260 12801
rect 24860 12656 24912 12708
rect 25780 12656 25832 12708
rect 29000 12656 29052 12708
rect 29092 12656 29144 12708
rect 30288 12724 30340 12776
rect 31392 12835 31444 12844
rect 31392 12801 31401 12835
rect 31401 12801 31435 12835
rect 31435 12801 31444 12835
rect 31392 12792 31444 12801
rect 25136 12631 25188 12640
rect 25136 12597 25145 12631
rect 25145 12597 25179 12631
rect 25179 12597 25188 12631
rect 25136 12588 25188 12597
rect 30012 12588 30064 12640
rect 31668 12724 31720 12776
rect 33876 12792 33928 12844
rect 32680 12724 32732 12776
rect 33324 12724 33376 12776
rect 32036 12656 32088 12708
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1676 12384 1728 12436
rect 3792 12427 3844 12436
rect 3792 12393 3801 12427
rect 3801 12393 3835 12427
rect 3835 12393 3844 12427
rect 3792 12384 3844 12393
rect 4068 12384 4120 12436
rect 4620 12384 4672 12436
rect 5816 12384 5868 12436
rect 8852 12384 8904 12436
rect 11152 12384 11204 12436
rect 16856 12427 16908 12436
rect 16856 12393 16865 12427
rect 16865 12393 16899 12427
rect 16899 12393 16908 12427
rect 16856 12384 16908 12393
rect 18328 12384 18380 12436
rect 19248 12384 19300 12436
rect 22376 12384 22428 12436
rect 3056 12291 3108 12300
rect 3056 12257 3065 12291
rect 3065 12257 3099 12291
rect 3099 12257 3108 12291
rect 3056 12248 3108 12257
rect 3240 12291 3292 12300
rect 3240 12257 3249 12291
rect 3249 12257 3283 12291
rect 3283 12257 3292 12291
rect 3240 12248 3292 12257
rect 4068 12248 4120 12300
rect 6276 12248 6328 12300
rect 7288 12248 7340 12300
rect 8852 12248 8904 12300
rect 3148 12112 3200 12164
rect 3424 12044 3476 12096
rect 8300 12180 8352 12232
rect 8760 12180 8812 12232
rect 10048 12180 10100 12232
rect 11980 12291 12032 12300
rect 11980 12257 11989 12291
rect 11989 12257 12023 12291
rect 12023 12257 12032 12291
rect 11980 12248 12032 12257
rect 12624 12248 12676 12300
rect 13176 12248 13228 12300
rect 16396 12316 16448 12368
rect 10232 12180 10284 12232
rect 14740 12223 14792 12232
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 14740 12180 14792 12189
rect 16488 12180 16540 12232
rect 7932 12112 7984 12164
rect 7840 12044 7892 12096
rect 9496 12112 9548 12164
rect 15292 12044 15344 12096
rect 17776 12248 17828 12300
rect 18328 12248 18380 12300
rect 19892 12316 19944 12368
rect 23572 12384 23624 12436
rect 18236 12180 18288 12232
rect 20812 12248 20864 12300
rect 23020 12291 23072 12300
rect 23020 12257 23029 12291
rect 23029 12257 23063 12291
rect 23063 12257 23072 12291
rect 23020 12248 23072 12257
rect 18972 12223 19024 12232
rect 18972 12189 18981 12223
rect 18981 12189 19015 12223
rect 19015 12189 19024 12223
rect 18972 12180 19024 12189
rect 19340 12223 19392 12232
rect 19340 12189 19349 12223
rect 19349 12189 19383 12223
rect 19383 12189 19392 12223
rect 19340 12180 19392 12189
rect 23296 12248 23348 12300
rect 24308 12384 24360 12436
rect 25136 12384 25188 12436
rect 25228 12427 25280 12436
rect 25228 12393 25237 12427
rect 25237 12393 25271 12427
rect 25271 12393 25280 12427
rect 25228 12384 25280 12393
rect 26332 12384 26384 12436
rect 26608 12384 26660 12436
rect 26792 12384 26844 12436
rect 29736 12384 29788 12436
rect 31760 12384 31812 12436
rect 32496 12384 32548 12436
rect 32680 12384 32732 12436
rect 32956 12384 33008 12436
rect 24768 12248 24820 12300
rect 26240 12291 26292 12300
rect 26240 12257 26249 12291
rect 26249 12257 26283 12291
rect 26283 12257 26292 12291
rect 26240 12248 26292 12257
rect 26332 12248 26384 12300
rect 27804 12248 27856 12300
rect 32312 12248 32364 12300
rect 20076 12112 20128 12164
rect 21456 12112 21508 12164
rect 23204 12223 23256 12232
rect 23204 12189 23213 12223
rect 23213 12189 23247 12223
rect 23247 12189 23256 12223
rect 23204 12180 23256 12189
rect 21824 12112 21876 12164
rect 23020 12112 23072 12164
rect 23848 12180 23900 12232
rect 24400 12180 24452 12232
rect 26424 12223 26476 12232
rect 26424 12189 26433 12223
rect 26433 12189 26467 12223
rect 26467 12189 26476 12223
rect 26424 12180 26476 12189
rect 27160 12180 27212 12232
rect 30012 12223 30064 12232
rect 30012 12189 30021 12223
rect 30021 12189 30055 12223
rect 30055 12189 30064 12223
rect 30012 12180 30064 12189
rect 17684 12044 17736 12096
rect 19432 12044 19484 12096
rect 22376 12044 22428 12096
rect 25780 12044 25832 12096
rect 26608 12044 26660 12096
rect 28448 12044 28500 12096
rect 28816 12044 28868 12096
rect 30472 12180 30524 12232
rect 33048 12180 33100 12232
rect 33232 12180 33284 12232
rect 30380 12044 30432 12096
rect 30472 12087 30524 12096
rect 30472 12053 30481 12087
rect 30481 12053 30515 12087
rect 30515 12053 30524 12087
rect 30472 12044 30524 12053
rect 32588 12044 32640 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 8760 11840 8812 11892
rect 9312 11840 9364 11892
rect 11336 11840 11388 11892
rect 12256 11840 12308 11892
rect 940 11704 992 11756
rect 8208 11704 8260 11756
rect 9312 11704 9364 11756
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 10324 11636 10376 11688
rect 10876 11679 10928 11688
rect 10876 11645 10885 11679
rect 10885 11645 10919 11679
rect 10919 11645 10928 11679
rect 10876 11636 10928 11645
rect 9588 11568 9640 11620
rect 14464 11840 14516 11892
rect 21272 11840 21324 11892
rect 22192 11840 22244 11892
rect 22652 11840 22704 11892
rect 27160 11840 27212 11892
rect 27620 11840 27672 11892
rect 29092 11840 29144 11892
rect 29368 11840 29420 11892
rect 30380 11840 30432 11892
rect 32680 11840 32732 11892
rect 15660 11772 15712 11824
rect 11888 11704 11940 11756
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 14832 11704 14884 11756
rect 12900 11636 12952 11688
rect 14280 11679 14332 11688
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 3608 11500 3660 11552
rect 8300 11500 8352 11552
rect 10324 11543 10376 11552
rect 10324 11509 10333 11543
rect 10333 11509 10367 11543
rect 10367 11509 10376 11543
rect 10324 11500 10376 11509
rect 15292 11636 15344 11688
rect 15568 11636 15620 11688
rect 18880 11772 18932 11824
rect 21824 11772 21876 11824
rect 22284 11772 22336 11824
rect 23572 11747 23624 11756
rect 23572 11713 23581 11747
rect 23581 11713 23615 11747
rect 23615 11713 23624 11747
rect 23572 11704 23624 11713
rect 24124 11704 24176 11756
rect 24216 11747 24268 11756
rect 24216 11713 24225 11747
rect 24225 11713 24259 11747
rect 24259 11713 24268 11747
rect 24216 11704 24268 11713
rect 24400 11704 24452 11756
rect 23480 11636 23532 11688
rect 23940 11636 23992 11688
rect 17592 11568 17644 11620
rect 18696 11611 18748 11620
rect 18696 11577 18705 11611
rect 18705 11577 18739 11611
rect 18739 11577 18748 11611
rect 18696 11568 18748 11577
rect 22100 11568 22152 11620
rect 24676 11704 24728 11756
rect 24768 11747 24820 11756
rect 24768 11713 24777 11747
rect 24777 11713 24811 11747
rect 24811 11713 24820 11747
rect 24768 11704 24820 11713
rect 26608 11772 26660 11824
rect 25044 11747 25096 11756
rect 25044 11713 25053 11747
rect 25053 11713 25087 11747
rect 25087 11713 25096 11747
rect 25044 11704 25096 11713
rect 26424 11636 26476 11688
rect 27436 11772 27488 11824
rect 27344 11747 27396 11756
rect 27344 11713 27353 11747
rect 27353 11713 27387 11747
rect 27387 11713 27396 11747
rect 27344 11704 27396 11713
rect 27804 11772 27856 11824
rect 27988 11772 28040 11824
rect 32220 11772 32272 11824
rect 28816 11704 28868 11756
rect 29000 11704 29052 11756
rect 29736 11704 29788 11756
rect 30288 11704 30340 11756
rect 30472 11704 30524 11756
rect 32588 11747 32640 11756
rect 32588 11713 32597 11747
rect 32597 11713 32631 11747
rect 32631 11713 32640 11747
rect 32588 11704 32640 11713
rect 33692 11704 33744 11756
rect 29828 11679 29880 11688
rect 29828 11645 29837 11679
rect 29837 11645 29871 11679
rect 29871 11645 29880 11679
rect 29828 11636 29880 11645
rect 30656 11679 30708 11688
rect 30656 11645 30665 11679
rect 30665 11645 30699 11679
rect 30699 11645 30708 11679
rect 30656 11636 30708 11645
rect 27160 11568 27212 11620
rect 27528 11611 27580 11620
rect 27528 11577 27537 11611
rect 27537 11577 27571 11611
rect 27571 11577 27580 11611
rect 27528 11568 27580 11577
rect 27896 11568 27948 11620
rect 34612 11568 34664 11620
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 19248 11500 19300 11552
rect 23480 11500 23532 11552
rect 25780 11500 25832 11552
rect 26884 11500 26936 11552
rect 27436 11500 27488 11552
rect 27712 11543 27764 11552
rect 27712 11509 27721 11543
rect 27721 11509 27755 11543
rect 27755 11509 27764 11543
rect 27712 11500 27764 11509
rect 27988 11500 28040 11552
rect 30288 11500 30340 11552
rect 30380 11500 30432 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3148 11339 3200 11348
rect 3148 11305 3157 11339
rect 3157 11305 3191 11339
rect 3191 11305 3200 11339
rect 3148 11296 3200 11305
rect 3424 11296 3476 11348
rect 5724 11339 5776 11348
rect 5724 11305 5733 11339
rect 5733 11305 5767 11339
rect 5767 11305 5776 11339
rect 5724 11296 5776 11305
rect 7840 11296 7892 11348
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 9128 11296 9180 11348
rect 3884 11228 3936 11280
rect 4068 11160 4120 11212
rect 5632 11160 5684 11212
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 1676 11067 1728 11076
rect 1676 11033 1685 11067
rect 1685 11033 1719 11067
rect 1719 11033 1728 11067
rect 1676 11024 1728 11033
rect 2964 11024 3016 11076
rect 3884 11024 3936 11076
rect 5816 11024 5868 11076
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 8208 11160 8260 11212
rect 8852 11228 8904 11280
rect 9312 11271 9364 11280
rect 9312 11237 9321 11271
rect 9321 11237 9355 11271
rect 9355 11237 9364 11271
rect 9312 11228 9364 11237
rect 9588 11228 9640 11280
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 8576 11092 8628 11101
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 10324 11296 10376 11348
rect 11980 11296 12032 11348
rect 14464 11296 14516 11348
rect 17592 11339 17644 11348
rect 17592 11305 17601 11339
rect 17601 11305 17635 11339
rect 17635 11305 17644 11339
rect 17592 11296 17644 11305
rect 19432 11296 19484 11348
rect 23480 11296 23532 11348
rect 25044 11296 25096 11348
rect 29184 11296 29236 11348
rect 30104 11296 30156 11348
rect 30380 11296 30432 11348
rect 30656 11296 30708 11348
rect 32128 11339 32180 11348
rect 32128 11305 32137 11339
rect 32137 11305 32171 11339
rect 32171 11305 32180 11339
rect 32128 11296 32180 11305
rect 32680 11296 32732 11348
rect 34612 11296 34664 11348
rect 9864 11160 9916 11212
rect 10784 11160 10836 11212
rect 12900 11203 12952 11212
rect 12900 11169 12909 11203
rect 12909 11169 12943 11203
rect 12943 11169 12952 11203
rect 12900 11160 12952 11169
rect 12624 11092 12676 11144
rect 7564 11024 7616 11076
rect 7840 11024 7892 11076
rect 8116 11024 8168 11076
rect 11336 11024 11388 11076
rect 12808 11067 12860 11076
rect 12808 11033 12817 11067
rect 12817 11033 12851 11067
rect 12851 11033 12860 11067
rect 12808 11024 12860 11033
rect 13360 11024 13412 11076
rect 15292 11228 15344 11280
rect 14832 11160 14884 11212
rect 18788 11228 18840 11280
rect 19248 11228 19300 11280
rect 15568 11135 15620 11144
rect 15568 11101 15577 11135
rect 15577 11101 15611 11135
rect 15611 11101 15620 11135
rect 15568 11092 15620 11101
rect 15752 11092 15804 11144
rect 18236 11092 18288 11144
rect 20260 11228 20312 11280
rect 21824 11228 21876 11280
rect 22284 11228 22336 11280
rect 23572 11228 23624 11280
rect 20076 11135 20128 11144
rect 20076 11101 20085 11135
rect 20085 11101 20119 11135
rect 20119 11101 20128 11135
rect 20076 11092 20128 11101
rect 22376 11160 22428 11212
rect 23112 11160 23164 11212
rect 26608 11228 26660 11280
rect 27068 11228 27120 11280
rect 20996 11024 21048 11076
rect 23664 11092 23716 11144
rect 3792 10999 3844 11008
rect 3792 10965 3801 10999
rect 3801 10965 3835 10999
rect 3835 10965 3844 10999
rect 3792 10956 3844 10965
rect 4252 10999 4304 11008
rect 4252 10965 4261 10999
rect 4261 10965 4295 10999
rect 4295 10965 4304 10999
rect 4252 10956 4304 10965
rect 6736 10956 6788 11008
rect 12348 10956 12400 11008
rect 14096 10956 14148 11008
rect 15936 10956 15988 11008
rect 16488 10956 16540 11008
rect 17040 10956 17092 11008
rect 21456 10956 21508 11008
rect 22100 11024 22152 11076
rect 21824 10956 21876 11008
rect 23296 11024 23348 11076
rect 24216 11160 24268 11212
rect 24768 11160 24820 11212
rect 26332 11160 26384 11212
rect 26240 11092 26292 11144
rect 26424 11135 26476 11144
rect 26424 11101 26433 11135
rect 26433 11101 26467 11135
rect 26467 11101 26476 11135
rect 26424 11092 26476 11101
rect 26516 11092 26568 11144
rect 27068 11135 27120 11144
rect 27068 11101 27077 11135
rect 27077 11101 27111 11135
rect 27111 11101 27120 11135
rect 27068 11092 27120 11101
rect 27344 11228 27396 11280
rect 27436 11228 27488 11280
rect 27620 11160 27672 11212
rect 27804 11092 27856 11144
rect 27988 11092 28040 11144
rect 31760 11228 31812 11280
rect 30472 11160 30524 11212
rect 29644 11092 29696 11144
rect 30196 11135 30248 11144
rect 30196 11101 30205 11135
rect 30205 11101 30239 11135
rect 30239 11101 30248 11135
rect 30196 11092 30248 11101
rect 30288 11135 30340 11144
rect 30288 11101 30297 11135
rect 30297 11101 30331 11135
rect 30331 11101 30340 11135
rect 30288 11092 30340 11101
rect 31852 11135 31904 11144
rect 31852 11101 31861 11135
rect 31861 11101 31895 11135
rect 31895 11101 31904 11135
rect 31852 11092 31904 11101
rect 32312 11135 32364 11144
rect 32312 11101 32321 11135
rect 32321 11101 32355 11135
rect 32355 11101 32364 11135
rect 32312 11092 32364 11101
rect 32496 11092 32548 11144
rect 32772 11135 32824 11144
rect 32772 11101 32781 11135
rect 32781 11101 32815 11135
rect 32815 11101 32824 11135
rect 32772 11092 32824 11101
rect 23388 10999 23440 11008
rect 23388 10965 23397 10999
rect 23397 10965 23431 10999
rect 23431 10965 23440 10999
rect 23388 10956 23440 10965
rect 25780 10956 25832 11008
rect 26792 10999 26844 11008
rect 26792 10965 26801 10999
rect 26801 10965 26835 10999
rect 26835 10965 26844 10999
rect 26792 10956 26844 10965
rect 27068 10956 27120 11008
rect 27620 10999 27672 11008
rect 27620 10965 27629 10999
rect 27629 10965 27663 10999
rect 27663 10965 27672 10999
rect 27620 10956 27672 10965
rect 30196 10956 30248 11008
rect 30656 10956 30708 11008
rect 37924 11067 37976 11076
rect 37924 11033 37933 11067
rect 37933 11033 37967 11067
rect 37967 11033 37976 11067
rect 37924 11024 37976 11033
rect 32588 10956 32640 11008
rect 32956 10999 33008 11008
rect 32956 10965 32965 10999
rect 32965 10965 32999 10999
rect 32999 10965 33008 10999
rect 32956 10956 33008 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1676 10752 1728 10804
rect 3792 10752 3844 10804
rect 3884 10752 3936 10804
rect 3148 10616 3200 10668
rect 3424 10591 3476 10600
rect 3424 10557 3433 10591
rect 3433 10557 3467 10591
rect 3467 10557 3476 10591
rect 3424 10548 3476 10557
rect 4252 10684 4304 10736
rect 6092 10752 6144 10804
rect 5632 10684 5684 10736
rect 8484 10752 8536 10804
rect 9404 10752 9456 10804
rect 5724 10616 5776 10668
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 4712 10548 4764 10600
rect 5816 10548 5868 10600
rect 15752 10752 15804 10804
rect 18880 10752 18932 10804
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7196 10616 7248 10625
rect 7472 10616 7524 10668
rect 8484 10616 8536 10668
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 10784 10616 10836 10668
rect 3240 10412 3292 10464
rect 5816 10412 5868 10464
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 8300 10412 8352 10464
rect 10232 10548 10284 10600
rect 11244 10591 11296 10600
rect 11244 10557 11253 10591
rect 11253 10557 11287 10591
rect 11287 10557 11296 10591
rect 11244 10548 11296 10557
rect 14096 10684 14148 10736
rect 15936 10727 15988 10736
rect 15936 10693 15945 10727
rect 15945 10693 15979 10727
rect 15979 10693 15988 10727
rect 15936 10684 15988 10693
rect 21548 10752 21600 10804
rect 15292 10616 15344 10668
rect 16488 10616 16540 10668
rect 16948 10616 17000 10668
rect 12256 10548 12308 10600
rect 17132 10659 17184 10668
rect 17132 10625 17141 10659
rect 17141 10625 17175 10659
rect 17175 10625 17184 10659
rect 17132 10616 17184 10625
rect 17500 10523 17552 10532
rect 17500 10489 17509 10523
rect 17509 10489 17543 10523
rect 17543 10489 17552 10523
rect 17500 10480 17552 10489
rect 18236 10616 18288 10668
rect 18788 10616 18840 10668
rect 20996 10727 21048 10736
rect 20996 10693 21021 10727
rect 21021 10693 21048 10727
rect 20996 10684 21048 10693
rect 22928 10684 22980 10736
rect 23112 10727 23164 10736
rect 23112 10693 23121 10727
rect 23121 10693 23155 10727
rect 23155 10693 23164 10727
rect 23112 10684 23164 10693
rect 23388 10684 23440 10736
rect 21180 10548 21232 10600
rect 21640 10591 21692 10600
rect 21640 10557 21649 10591
rect 21649 10557 21683 10591
rect 21683 10557 21692 10591
rect 21640 10548 21692 10557
rect 21916 10591 21968 10600
rect 21916 10557 21925 10591
rect 21925 10557 21959 10591
rect 21959 10557 21968 10591
rect 22376 10659 22428 10668
rect 22376 10625 22385 10659
rect 22385 10625 22419 10659
rect 22419 10625 22428 10659
rect 22376 10616 22428 10625
rect 22468 10659 22520 10668
rect 22468 10625 22477 10659
rect 22477 10625 22511 10659
rect 22511 10625 22520 10659
rect 22468 10616 22520 10625
rect 22836 10616 22888 10668
rect 21916 10548 21968 10557
rect 20812 10480 20864 10532
rect 21824 10480 21876 10532
rect 23112 10548 23164 10600
rect 23296 10548 23348 10600
rect 23480 10616 23532 10668
rect 24400 10752 24452 10804
rect 27620 10752 27672 10804
rect 28172 10752 28224 10804
rect 26792 10616 26844 10668
rect 27252 10659 27304 10668
rect 27252 10625 27261 10659
rect 27261 10625 27295 10659
rect 27295 10625 27304 10659
rect 27252 10616 27304 10625
rect 27528 10616 27580 10668
rect 28448 10684 28500 10736
rect 32312 10752 32364 10804
rect 32588 10752 32640 10804
rect 33692 10795 33744 10804
rect 33692 10761 33701 10795
rect 33701 10761 33735 10795
rect 33735 10761 33744 10795
rect 33692 10752 33744 10761
rect 35624 10752 35676 10804
rect 29092 10684 29144 10736
rect 28356 10659 28408 10668
rect 28356 10625 28365 10659
rect 28365 10625 28399 10659
rect 28399 10625 28408 10659
rect 28356 10616 28408 10625
rect 28816 10616 28868 10668
rect 29000 10616 29052 10668
rect 30288 10659 30340 10668
rect 30288 10625 30297 10659
rect 30297 10625 30331 10659
rect 30331 10625 30340 10659
rect 30288 10616 30340 10625
rect 31852 10616 31904 10668
rect 32220 10616 32272 10668
rect 32772 10616 32824 10668
rect 33508 10659 33560 10668
rect 33508 10625 33517 10659
rect 33517 10625 33551 10659
rect 33551 10625 33560 10659
rect 33508 10616 33560 10625
rect 23756 10548 23808 10600
rect 24400 10548 24452 10600
rect 17040 10412 17092 10464
rect 18052 10455 18104 10464
rect 18052 10421 18061 10455
rect 18061 10421 18095 10455
rect 18095 10421 18104 10455
rect 18052 10412 18104 10421
rect 20168 10455 20220 10464
rect 20168 10421 20177 10455
rect 20177 10421 20211 10455
rect 20211 10421 20220 10455
rect 20168 10412 20220 10421
rect 21088 10412 21140 10464
rect 21640 10412 21692 10464
rect 22376 10412 22428 10464
rect 22744 10455 22796 10464
rect 22744 10421 22753 10455
rect 22753 10421 22787 10455
rect 22787 10421 22796 10455
rect 22744 10412 22796 10421
rect 24032 10412 24084 10464
rect 28172 10480 28224 10532
rect 32496 10591 32548 10600
rect 32496 10557 32505 10591
rect 32505 10557 32539 10591
rect 32539 10557 32548 10591
rect 32496 10548 32548 10557
rect 33232 10548 33284 10600
rect 27896 10412 27948 10464
rect 32128 10412 32180 10464
rect 32864 10455 32916 10464
rect 32864 10421 32873 10455
rect 32873 10421 32907 10455
rect 32907 10421 32916 10455
rect 32864 10412 32916 10421
rect 34428 10616 34480 10668
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4712 10208 4764 10260
rect 6184 10251 6236 10260
rect 6184 10217 6193 10251
rect 6193 10217 6227 10251
rect 6227 10217 6236 10251
rect 6184 10208 6236 10217
rect 6368 10208 6420 10260
rect 7564 10251 7616 10260
rect 7564 10217 7573 10251
rect 7573 10217 7607 10251
rect 7607 10217 7616 10251
rect 7564 10208 7616 10217
rect 9956 10208 10008 10260
rect 11796 10208 11848 10260
rect 12164 10208 12216 10260
rect 12348 10208 12400 10260
rect 13084 10208 13136 10260
rect 13912 10208 13964 10260
rect 14372 10208 14424 10260
rect 17132 10208 17184 10260
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 5908 10072 5960 10124
rect 3148 10004 3200 10056
rect 3332 10004 3384 10056
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 6092 10004 6144 10056
rect 7472 10047 7524 10056
rect 7472 10013 7481 10047
rect 7481 10013 7515 10047
rect 7515 10013 7524 10047
rect 7472 10004 7524 10013
rect 8024 10140 8076 10192
rect 8208 10072 8260 10124
rect 8668 10072 8720 10124
rect 7932 10004 7984 10056
rect 8944 10004 8996 10056
rect 9496 10140 9548 10192
rect 10692 10140 10744 10192
rect 9772 10072 9824 10124
rect 18696 10208 18748 10260
rect 19248 10208 19300 10260
rect 20260 10208 20312 10260
rect 20536 10140 20588 10192
rect 8484 9936 8536 9988
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 13268 10004 13320 10056
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 9496 9911 9548 9920
rect 9496 9877 9505 9911
rect 9505 9877 9539 9911
rect 9539 9877 9548 9911
rect 9496 9868 9548 9877
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 18236 10047 18288 10056
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 18328 10047 18380 10056
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 18788 10004 18840 10056
rect 20168 10004 20220 10056
rect 20444 10047 20496 10056
rect 20444 10013 20453 10047
rect 20453 10013 20487 10047
rect 20487 10013 20496 10047
rect 20444 10004 20496 10013
rect 21824 10208 21876 10260
rect 22376 10251 22428 10260
rect 22376 10217 22385 10251
rect 22385 10217 22419 10251
rect 22419 10217 22428 10251
rect 22376 10208 22428 10217
rect 22468 10208 22520 10260
rect 22744 10208 22796 10260
rect 25688 10208 25740 10260
rect 28448 10208 28500 10260
rect 12164 9868 12216 9920
rect 20352 9936 20404 9988
rect 20628 9979 20680 9988
rect 20628 9945 20637 9979
rect 20637 9945 20671 9979
rect 20671 9945 20680 9979
rect 20628 9936 20680 9945
rect 20904 9936 20956 9988
rect 21180 10004 21232 10056
rect 24124 10140 24176 10192
rect 28908 10140 28960 10192
rect 29092 10140 29144 10192
rect 30748 10208 30800 10260
rect 32772 10208 32824 10260
rect 33508 10251 33560 10260
rect 33508 10217 33517 10251
rect 33517 10217 33551 10251
rect 33551 10217 33560 10251
rect 33508 10208 33560 10217
rect 26424 10072 26476 10124
rect 27896 10072 27948 10124
rect 28172 10072 28224 10124
rect 21640 10047 21692 10056
rect 21640 10013 21649 10047
rect 21649 10013 21683 10047
rect 21683 10013 21692 10047
rect 21640 10004 21692 10013
rect 21824 10047 21876 10056
rect 21824 10013 21833 10047
rect 21833 10013 21867 10047
rect 21867 10013 21876 10047
rect 21824 10004 21876 10013
rect 22192 10004 22244 10056
rect 22284 10047 22336 10056
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 22560 10004 22612 10056
rect 26148 10004 26200 10056
rect 28356 10004 28408 10056
rect 28724 10047 28776 10056
rect 28724 10013 28733 10047
rect 28733 10013 28767 10047
rect 28767 10013 28776 10047
rect 28724 10004 28776 10013
rect 28908 10047 28960 10056
rect 28908 10013 28917 10047
rect 28917 10013 28951 10047
rect 28951 10013 28960 10047
rect 28908 10004 28960 10013
rect 30380 10115 30432 10124
rect 30380 10081 30389 10115
rect 30389 10081 30423 10115
rect 30423 10081 30432 10115
rect 30380 10072 30432 10081
rect 30196 10004 30248 10056
rect 30656 10047 30708 10056
rect 30656 10013 30665 10047
rect 30665 10013 30699 10047
rect 30699 10013 30708 10047
rect 32956 10140 33008 10192
rect 30656 10004 30708 10013
rect 32864 10004 32916 10056
rect 13452 9868 13504 9920
rect 16672 9868 16724 9920
rect 26332 9936 26384 9988
rect 27896 9936 27948 9988
rect 29000 9936 29052 9988
rect 33968 10047 34020 10056
rect 33968 10013 33977 10047
rect 33977 10013 34011 10047
rect 34011 10013 34020 10047
rect 33968 10004 34020 10013
rect 34060 10004 34112 10056
rect 22928 9868 22980 9920
rect 24860 9868 24912 9920
rect 24952 9868 25004 9920
rect 28908 9868 28960 9920
rect 30840 9911 30892 9920
rect 30840 9877 30849 9911
rect 30849 9877 30883 9911
rect 30883 9877 30892 9911
rect 30840 9868 30892 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 3148 9664 3200 9716
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 5540 9596 5592 9648
rect 8208 9596 8260 9648
rect 11428 9664 11480 9716
rect 13084 9707 13136 9716
rect 13084 9673 13093 9707
rect 13093 9673 13127 9707
rect 13127 9673 13136 9707
rect 13084 9664 13136 9673
rect 13452 9707 13504 9716
rect 13452 9673 13461 9707
rect 13461 9673 13495 9707
rect 13495 9673 13504 9707
rect 13452 9664 13504 9673
rect 10600 9596 10652 9648
rect 11612 9596 11664 9648
rect 11704 9596 11756 9648
rect 13176 9596 13228 9648
rect 3700 9528 3752 9580
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 7104 9528 7156 9580
rect 7840 9528 7892 9580
rect 8116 9528 8168 9580
rect 8484 9571 8536 9580
rect 8484 9537 8493 9571
rect 8493 9537 8527 9571
rect 8527 9537 8536 9571
rect 8484 9528 8536 9537
rect 8944 9528 8996 9580
rect 7472 9435 7524 9444
rect 7472 9401 7481 9435
rect 7481 9401 7515 9435
rect 7515 9401 7524 9435
rect 7472 9392 7524 9401
rect 8208 9392 8260 9444
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 14372 9596 14424 9648
rect 13728 9528 13780 9580
rect 13820 9528 13872 9580
rect 14096 9528 14148 9580
rect 15292 9596 15344 9648
rect 15384 9528 15436 9580
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 12624 9460 12676 9512
rect 13268 9460 13320 9512
rect 15200 9460 15252 9512
rect 15660 9460 15712 9512
rect 20260 9664 20312 9716
rect 22376 9664 22428 9716
rect 18052 9596 18104 9648
rect 16672 9528 16724 9580
rect 17316 9528 17368 9580
rect 18328 9528 18380 9580
rect 19892 9571 19944 9580
rect 19892 9537 19901 9571
rect 19901 9537 19935 9571
rect 19935 9537 19944 9571
rect 19892 9528 19944 9537
rect 20168 9528 20220 9580
rect 23020 9664 23072 9716
rect 23480 9664 23532 9716
rect 23572 9664 23624 9716
rect 23756 9596 23808 9648
rect 24124 9664 24176 9716
rect 24860 9664 24912 9716
rect 27344 9664 27396 9716
rect 16948 9460 17000 9512
rect 17500 9460 17552 9512
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 3976 9324 4028 9376
rect 4712 9324 4764 9376
rect 7288 9324 7340 9376
rect 9680 9324 9732 9376
rect 10048 9367 10100 9376
rect 10048 9333 10057 9367
rect 10057 9333 10091 9367
rect 10091 9333 10100 9367
rect 10048 9324 10100 9333
rect 11428 9392 11480 9444
rect 12164 9392 12216 9444
rect 18328 9392 18380 9444
rect 13176 9324 13228 9376
rect 13912 9324 13964 9376
rect 16028 9367 16080 9376
rect 16028 9333 16037 9367
rect 16037 9333 16071 9367
rect 16071 9333 16080 9367
rect 16028 9324 16080 9333
rect 16304 9324 16356 9376
rect 19432 9503 19484 9512
rect 19432 9469 19441 9503
rect 19441 9469 19475 9503
rect 19475 9469 19484 9503
rect 19432 9460 19484 9469
rect 20260 9460 20312 9512
rect 19064 9392 19116 9444
rect 22284 9392 22336 9444
rect 22744 9392 22796 9444
rect 19340 9324 19392 9376
rect 22560 9324 22612 9376
rect 23388 9528 23440 9580
rect 24952 9596 25004 9648
rect 33140 9664 33192 9716
rect 33968 9664 34020 9716
rect 23296 9460 23348 9512
rect 25504 9460 25556 9512
rect 26148 9571 26200 9580
rect 26148 9537 26157 9571
rect 26157 9537 26191 9571
rect 26191 9537 26200 9571
rect 26148 9528 26200 9537
rect 27068 9528 27120 9580
rect 27344 9528 27396 9580
rect 24308 9435 24360 9444
rect 24308 9401 24317 9435
rect 24317 9401 24351 9435
rect 24351 9401 24360 9435
rect 24308 9392 24360 9401
rect 27712 9528 27764 9580
rect 28724 9528 28776 9580
rect 28908 9528 28960 9580
rect 29644 9571 29696 9580
rect 29644 9537 29653 9571
rect 29653 9537 29687 9571
rect 29687 9537 29696 9571
rect 29644 9528 29696 9537
rect 29736 9571 29788 9580
rect 29736 9537 29745 9571
rect 29745 9537 29779 9571
rect 29779 9537 29788 9571
rect 29736 9528 29788 9537
rect 30104 9571 30156 9580
rect 30104 9537 30113 9571
rect 30113 9537 30147 9571
rect 30147 9537 30156 9571
rect 30104 9528 30156 9537
rect 30748 9571 30800 9580
rect 30748 9537 30757 9571
rect 30757 9537 30791 9571
rect 30791 9537 30800 9571
rect 30748 9528 30800 9537
rect 30840 9528 30892 9580
rect 31392 9528 31444 9580
rect 30196 9460 30248 9512
rect 24124 9324 24176 9376
rect 26516 9367 26568 9376
rect 26516 9333 26525 9367
rect 26525 9333 26559 9367
rect 26559 9333 26568 9367
rect 30932 9392 30984 9444
rect 33048 9639 33100 9648
rect 33048 9605 33057 9639
rect 33057 9605 33091 9639
rect 33091 9605 33100 9639
rect 33048 9596 33100 9605
rect 32772 9528 32824 9580
rect 32036 9392 32088 9444
rect 26516 9324 26568 9333
rect 28080 9324 28132 9376
rect 29736 9324 29788 9376
rect 31576 9324 31628 9376
rect 31668 9324 31720 9376
rect 33232 9324 33284 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2964 9120 3016 9172
rect 6828 9120 6880 9172
rect 7104 9120 7156 9172
rect 3976 9052 4028 9104
rect 3332 8916 3384 8968
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 6736 9052 6788 9104
rect 4712 8984 4764 9036
rect 11612 9120 11664 9172
rect 14096 9120 14148 9172
rect 15292 9120 15344 9172
rect 18236 9120 18288 9172
rect 18328 9120 18380 9172
rect 19064 9120 19116 9172
rect 21088 9120 21140 9172
rect 22100 9120 22152 9172
rect 940 8848 992 8900
rect 3884 8823 3936 8832
rect 3884 8789 3893 8823
rect 3893 8789 3927 8823
rect 3927 8789 3936 8823
rect 3884 8780 3936 8789
rect 4712 8848 4764 8900
rect 7196 8916 7248 8968
rect 6000 8891 6052 8900
rect 6000 8857 6009 8891
rect 6009 8857 6043 8891
rect 6043 8857 6052 8891
rect 6000 8848 6052 8857
rect 5816 8780 5868 8832
rect 6184 8848 6236 8900
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 10600 8984 10652 9036
rect 11336 8916 11388 8968
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 13728 8984 13780 9036
rect 13820 8916 13872 8968
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 8484 8823 8536 8832
rect 8484 8789 8493 8823
rect 8493 8789 8527 8823
rect 8527 8789 8536 8823
rect 8484 8780 8536 8789
rect 9956 8848 10008 8900
rect 11428 8848 11480 8900
rect 11704 8848 11756 8900
rect 14372 8959 14424 8968
rect 14372 8925 14384 8959
rect 14384 8925 14418 8959
rect 14418 8925 14424 8959
rect 14372 8916 14424 8925
rect 15016 8916 15068 8968
rect 18972 9052 19024 9104
rect 15384 8984 15436 9036
rect 17592 8984 17644 9036
rect 20260 9027 20312 9036
rect 15752 8959 15804 8968
rect 15752 8925 15761 8959
rect 15761 8925 15795 8959
rect 15795 8925 15804 8959
rect 15752 8916 15804 8925
rect 15936 8848 15988 8900
rect 16028 8891 16080 8900
rect 16028 8857 16037 8891
rect 16037 8857 16071 8891
rect 16071 8857 16080 8891
rect 16028 8848 16080 8857
rect 16764 8848 16816 8900
rect 13084 8780 13136 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 14648 8780 14700 8832
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 14924 8823 14976 8832
rect 14924 8789 14933 8823
rect 14933 8789 14967 8823
rect 14967 8789 14976 8823
rect 14924 8780 14976 8789
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18696 8916 18748 8925
rect 20260 8993 20269 9027
rect 20269 8993 20303 9027
rect 20303 8993 20312 9027
rect 20260 8984 20312 8993
rect 20352 8984 20404 9036
rect 22192 9027 22244 9036
rect 22192 8993 22201 9027
rect 22201 8993 22235 9027
rect 22235 8993 22244 9027
rect 22192 8984 22244 8993
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 19984 8959 20036 8968
rect 19984 8925 19993 8959
rect 19993 8925 20027 8959
rect 20027 8925 20036 8959
rect 19984 8916 20036 8925
rect 20628 8959 20680 8968
rect 20628 8925 20637 8959
rect 20637 8925 20671 8959
rect 20671 8925 20680 8959
rect 20628 8916 20680 8925
rect 22560 8959 22612 8968
rect 22560 8925 22569 8959
rect 22569 8925 22603 8959
rect 22603 8925 22612 8959
rect 22560 8916 22612 8925
rect 20076 8848 20128 8900
rect 20168 8848 20220 8900
rect 22284 8891 22336 8900
rect 22284 8857 22293 8891
rect 22293 8857 22327 8891
rect 22327 8857 22336 8891
rect 22284 8848 22336 8857
rect 22928 9052 22980 9104
rect 23112 9052 23164 9104
rect 24400 9052 24452 9104
rect 24584 9052 24636 9104
rect 24860 9052 24912 9104
rect 26608 9120 26660 9172
rect 27252 9120 27304 9172
rect 29736 9163 29788 9172
rect 29736 9129 29745 9163
rect 29745 9129 29779 9163
rect 29779 9129 29788 9163
rect 29736 9120 29788 9129
rect 23020 8959 23072 8968
rect 23020 8925 23030 8959
rect 23030 8925 23064 8959
rect 23064 8925 23072 8959
rect 23020 8916 23072 8925
rect 23388 8959 23440 8968
rect 23388 8925 23402 8959
rect 23402 8925 23436 8959
rect 23436 8925 23440 8959
rect 23388 8916 23440 8925
rect 23756 8916 23808 8968
rect 24400 8959 24452 8968
rect 24400 8925 24409 8959
rect 24409 8925 24443 8959
rect 24443 8925 24452 8959
rect 24400 8916 24452 8925
rect 23296 8891 23348 8900
rect 23296 8857 23305 8891
rect 23305 8857 23339 8891
rect 23339 8857 23348 8891
rect 24952 8916 25004 8968
rect 23296 8848 23348 8857
rect 24584 8848 24636 8900
rect 20352 8780 20404 8832
rect 21824 8780 21876 8832
rect 23572 8823 23624 8832
rect 23572 8789 23581 8823
rect 23581 8789 23615 8823
rect 23615 8789 23624 8823
rect 23572 8780 23624 8789
rect 25136 8780 25188 8832
rect 25412 8916 25464 8968
rect 25872 8959 25924 8968
rect 25872 8925 25881 8959
rect 25881 8925 25915 8959
rect 25915 8925 25924 8959
rect 25872 8916 25924 8925
rect 27160 9052 27212 9104
rect 26516 8984 26568 9036
rect 25320 8848 25372 8900
rect 25780 8848 25832 8900
rect 26792 8959 26844 8968
rect 26792 8925 26801 8959
rect 26801 8925 26835 8959
rect 26835 8925 26844 8959
rect 26792 8916 26844 8925
rect 27804 8984 27856 9036
rect 28080 8984 28132 9036
rect 26976 8959 27028 8968
rect 26976 8925 26985 8959
rect 26985 8925 27019 8959
rect 27019 8925 27028 8959
rect 26976 8916 27028 8925
rect 27160 8959 27212 8968
rect 27160 8925 27169 8959
rect 27169 8925 27203 8959
rect 27203 8925 27212 8959
rect 27160 8916 27212 8925
rect 27252 8916 27304 8968
rect 27988 8959 28040 8968
rect 27988 8925 27997 8959
rect 27997 8925 28031 8959
rect 28031 8925 28040 8959
rect 27988 8916 28040 8925
rect 26332 8780 26384 8832
rect 26516 8823 26568 8832
rect 26516 8789 26525 8823
rect 26525 8789 26559 8823
rect 26559 8789 26568 8823
rect 26516 8780 26568 8789
rect 27712 8848 27764 8900
rect 28448 8959 28500 8968
rect 28448 8925 28457 8959
rect 28457 8925 28491 8959
rect 28491 8925 28500 8959
rect 28448 8916 28500 8925
rect 29184 9052 29236 9104
rect 29828 9052 29880 9104
rect 29368 8959 29420 8968
rect 29368 8925 29377 8959
rect 29377 8925 29411 8959
rect 29411 8925 29420 8959
rect 29368 8916 29420 8925
rect 29276 8848 29328 8900
rect 28816 8823 28868 8832
rect 28816 8789 28825 8823
rect 28825 8789 28859 8823
rect 28859 8789 28868 8823
rect 28816 8780 28868 8789
rect 28908 8780 28960 8832
rect 29000 8823 29052 8832
rect 29000 8789 29009 8823
rect 29009 8789 29043 8823
rect 29043 8789 29052 8823
rect 29000 8780 29052 8789
rect 29092 8780 29144 8832
rect 30104 8916 30156 8968
rect 30380 8891 30432 8900
rect 30380 8857 30389 8891
rect 30389 8857 30423 8891
rect 30423 8857 30432 8891
rect 30380 8848 30432 8857
rect 30748 9120 30800 9172
rect 31576 9120 31628 9172
rect 33140 9120 33192 9172
rect 33324 9120 33376 9172
rect 32036 8984 32088 9036
rect 31760 8916 31812 8968
rect 31852 8959 31904 8968
rect 31852 8925 31861 8959
rect 31861 8925 31895 8959
rect 31895 8925 31904 8959
rect 31852 8916 31904 8925
rect 30932 8780 30984 8832
rect 31944 8823 31996 8832
rect 31944 8789 31953 8823
rect 31953 8789 31987 8823
rect 31987 8789 31996 8823
rect 31944 8780 31996 8789
rect 32772 8916 32824 8968
rect 32864 8848 32916 8900
rect 33048 8959 33100 8968
rect 33048 8925 33057 8959
rect 33057 8925 33091 8959
rect 33091 8925 33100 8959
rect 33048 8916 33100 8925
rect 33140 8916 33192 8968
rect 38292 8916 38344 8968
rect 35900 8848 35952 8900
rect 36820 8848 36872 8900
rect 33232 8780 33284 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 5908 8576 5960 8628
rect 8484 8576 8536 8628
rect 10140 8576 10192 8628
rect 4712 8440 4764 8492
rect 4068 8304 4120 8356
rect 2964 8236 3016 8288
rect 4620 8236 4672 8288
rect 6000 8440 6052 8492
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 5632 8415 5684 8424
rect 5632 8381 5641 8415
rect 5641 8381 5675 8415
rect 5675 8381 5684 8415
rect 5632 8372 5684 8381
rect 6368 8440 6420 8492
rect 9404 8440 9456 8492
rect 9864 8440 9916 8492
rect 9956 8440 10008 8492
rect 11336 8576 11388 8628
rect 12256 8576 12308 8628
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 11152 8440 11204 8492
rect 11796 8440 11848 8492
rect 12624 8551 12676 8560
rect 12624 8517 12633 8551
rect 12633 8517 12667 8551
rect 12667 8517 12676 8551
rect 12624 8508 12676 8517
rect 13084 8508 13136 8560
rect 10416 8372 10468 8424
rect 11888 8415 11940 8424
rect 11888 8381 11897 8415
rect 11897 8381 11931 8415
rect 11931 8381 11940 8415
rect 11888 8372 11940 8381
rect 12164 8304 12216 8356
rect 5724 8236 5776 8288
rect 5908 8279 5960 8288
rect 5908 8245 5917 8279
rect 5917 8245 5951 8279
rect 5951 8245 5960 8279
rect 5908 8236 5960 8245
rect 6368 8236 6420 8288
rect 6828 8236 6880 8288
rect 8392 8236 8444 8288
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 14648 8576 14700 8628
rect 18420 8576 18472 8628
rect 18972 8576 19024 8628
rect 17316 8508 17368 8560
rect 20260 8576 20312 8628
rect 21824 8576 21876 8628
rect 16764 8440 16816 8492
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 18604 8440 18656 8492
rect 18880 8440 18932 8492
rect 18972 8483 19024 8492
rect 18972 8449 18981 8483
rect 18981 8449 19015 8483
rect 19015 8449 19024 8483
rect 18972 8440 19024 8449
rect 15016 8372 15068 8424
rect 19984 8440 20036 8492
rect 17224 8347 17276 8356
rect 17224 8313 17233 8347
rect 17233 8313 17267 8347
rect 17267 8313 17276 8347
rect 17224 8304 17276 8313
rect 20168 8372 20220 8424
rect 21640 8508 21692 8560
rect 22008 8440 22060 8492
rect 23572 8576 23624 8628
rect 24308 8576 24360 8628
rect 26976 8576 27028 8628
rect 28908 8576 28960 8628
rect 24124 8508 24176 8560
rect 23572 8440 23624 8492
rect 23848 8440 23900 8492
rect 24676 8440 24728 8492
rect 25320 8508 25372 8560
rect 26516 8440 26568 8492
rect 29000 8508 29052 8560
rect 30104 8576 30156 8628
rect 31392 8576 31444 8628
rect 32036 8576 32088 8628
rect 21916 8304 21968 8356
rect 23296 8372 23348 8424
rect 25412 8372 25464 8424
rect 26792 8372 26844 8424
rect 27068 8372 27120 8424
rect 27620 8440 27672 8492
rect 30196 8508 30248 8560
rect 31944 8508 31996 8560
rect 31668 8440 31720 8492
rect 29368 8372 29420 8424
rect 31024 8372 31076 8424
rect 35900 8508 35952 8560
rect 33048 8440 33100 8492
rect 12808 8236 12860 8288
rect 13728 8236 13780 8288
rect 15660 8236 15712 8288
rect 19524 8279 19576 8288
rect 19524 8245 19533 8279
rect 19533 8245 19567 8279
rect 19567 8245 19576 8279
rect 19524 8236 19576 8245
rect 22376 8236 22428 8288
rect 23020 8279 23072 8288
rect 23020 8245 23029 8279
rect 23029 8245 23063 8279
rect 23063 8245 23072 8279
rect 23020 8236 23072 8245
rect 25320 8279 25372 8288
rect 25320 8245 25329 8279
rect 25329 8245 25363 8279
rect 25363 8245 25372 8279
rect 25320 8236 25372 8245
rect 27528 8304 27580 8356
rect 27804 8304 27856 8356
rect 33232 8415 33284 8424
rect 33232 8381 33241 8415
rect 33241 8381 33275 8415
rect 33275 8381 33284 8415
rect 33232 8372 33284 8381
rect 32588 8304 32640 8356
rect 29000 8279 29052 8288
rect 29000 8245 29009 8279
rect 29009 8245 29043 8279
rect 29043 8245 29052 8279
rect 29000 8236 29052 8245
rect 29644 8236 29696 8288
rect 34060 8236 34112 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 5540 8032 5592 8084
rect 5816 8032 5868 8084
rect 5724 7828 5776 7880
rect 5908 7828 5960 7880
rect 8392 8032 8444 8084
rect 10508 8032 10560 8084
rect 11520 8032 11572 8084
rect 12256 8032 12308 8084
rect 12532 8032 12584 8084
rect 12992 8032 13044 8084
rect 13728 8075 13780 8084
rect 13728 8041 13737 8075
rect 13737 8041 13771 8075
rect 13771 8041 13780 8075
rect 13728 8032 13780 8041
rect 19432 8032 19484 8084
rect 23572 8032 23624 8084
rect 26240 8032 26292 8084
rect 29276 8032 29328 8084
rect 30840 8032 30892 8084
rect 31484 8032 31536 8084
rect 31760 8032 31812 8084
rect 20260 7964 20312 8016
rect 22652 7964 22704 8016
rect 22744 7964 22796 8016
rect 24032 7964 24084 8016
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 9404 7896 9456 7948
rect 9680 7871 9732 7880
rect 9680 7837 9697 7871
rect 9697 7837 9731 7871
rect 9731 7837 9732 7871
rect 11888 7896 11940 7948
rect 9680 7828 9732 7837
rect 7196 7803 7248 7812
rect 7196 7769 7205 7803
rect 7205 7769 7239 7803
rect 7239 7769 7248 7803
rect 7196 7760 7248 7769
rect 8484 7760 8536 7812
rect 9772 7760 9824 7812
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 9680 7735 9732 7744
rect 9680 7701 9689 7735
rect 9689 7701 9723 7735
rect 9723 7701 9732 7735
rect 9680 7692 9732 7701
rect 9956 7828 10008 7880
rect 10968 7828 11020 7880
rect 12348 7803 12400 7812
rect 12348 7769 12357 7803
rect 12357 7769 12391 7803
rect 12391 7769 12400 7803
rect 12348 7760 12400 7769
rect 10876 7692 10928 7744
rect 13636 7896 13688 7948
rect 14004 7896 14056 7948
rect 15660 7896 15712 7948
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 19524 7896 19576 7948
rect 17592 7871 17644 7880
rect 13636 7760 13688 7812
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 17776 7871 17828 7880
rect 17776 7837 17785 7871
rect 17785 7837 17819 7871
rect 17819 7837 17828 7871
rect 17776 7828 17828 7837
rect 20628 7896 20680 7948
rect 16856 7760 16908 7812
rect 21640 7828 21692 7880
rect 22284 7896 22336 7948
rect 22376 7939 22428 7948
rect 22376 7905 22385 7939
rect 22385 7905 22419 7939
rect 22419 7905 22428 7939
rect 22376 7896 22428 7905
rect 21824 7871 21876 7880
rect 21824 7837 21833 7871
rect 21833 7837 21867 7871
rect 21867 7837 21876 7871
rect 21824 7828 21876 7837
rect 23020 7896 23072 7948
rect 29000 7896 29052 7948
rect 29920 7896 29972 7948
rect 15384 7735 15436 7744
rect 15384 7701 15393 7735
rect 15393 7701 15427 7735
rect 15427 7701 15436 7735
rect 15384 7692 15436 7701
rect 17316 7735 17368 7744
rect 17316 7701 17325 7735
rect 17325 7701 17359 7735
rect 17359 7701 17368 7735
rect 17316 7692 17368 7701
rect 20536 7692 20588 7744
rect 22652 7871 22704 7880
rect 22652 7837 22661 7871
rect 22661 7837 22695 7871
rect 22695 7837 22704 7871
rect 22652 7828 22704 7837
rect 30012 7871 30064 7880
rect 30012 7837 30021 7871
rect 30021 7837 30055 7871
rect 30055 7837 30064 7871
rect 30012 7828 30064 7837
rect 30472 7896 30524 7948
rect 33048 7964 33100 8016
rect 31116 7896 31168 7948
rect 30380 7871 30432 7880
rect 30380 7837 30389 7871
rect 30389 7837 30423 7871
rect 30423 7837 30432 7871
rect 30380 7828 30432 7837
rect 22376 7760 22428 7812
rect 22560 7760 22612 7812
rect 23112 7803 23164 7812
rect 23112 7769 23121 7803
rect 23121 7769 23155 7803
rect 23155 7769 23164 7803
rect 23112 7760 23164 7769
rect 25044 7760 25096 7812
rect 25872 7760 25924 7812
rect 27344 7760 27396 7812
rect 30840 7828 30892 7880
rect 30932 7871 30984 7880
rect 30932 7837 30941 7871
rect 30941 7837 30975 7871
rect 30975 7837 30984 7871
rect 30932 7828 30984 7837
rect 31024 7828 31076 7880
rect 31668 7803 31720 7812
rect 31668 7769 31677 7803
rect 31677 7769 31711 7803
rect 31711 7769 31720 7803
rect 31668 7760 31720 7769
rect 22100 7692 22152 7744
rect 22284 7735 22336 7744
rect 22284 7701 22293 7735
rect 22293 7701 22327 7735
rect 22327 7701 22336 7735
rect 22284 7692 22336 7701
rect 30564 7692 30616 7744
rect 31208 7735 31260 7744
rect 31208 7701 31217 7735
rect 31217 7701 31251 7735
rect 31251 7701 31260 7735
rect 31208 7692 31260 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 4620 7488 4672 7540
rect 6092 7488 6144 7540
rect 6552 7488 6604 7540
rect 7196 7488 7248 7540
rect 8024 7488 8076 7540
rect 13176 7488 13228 7540
rect 2964 7420 3016 7472
rect 3976 7352 4028 7404
rect 6000 7352 6052 7404
rect 3608 7284 3660 7336
rect 4712 7284 4764 7336
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 9772 7420 9824 7472
rect 11796 7463 11848 7472
rect 11796 7429 11805 7463
rect 11805 7429 11839 7463
rect 11839 7429 11848 7463
rect 11796 7420 11848 7429
rect 12440 7420 12492 7472
rect 14648 7420 14700 7472
rect 15384 7488 15436 7540
rect 18604 7488 18656 7540
rect 15292 7352 15344 7404
rect 21364 7488 21416 7540
rect 22284 7488 22336 7540
rect 22376 7531 22428 7540
rect 22376 7497 22385 7531
rect 22385 7497 22419 7531
rect 22419 7497 22428 7531
rect 22376 7488 22428 7497
rect 17776 7395 17828 7404
rect 17776 7361 17785 7395
rect 17785 7361 17819 7395
rect 17819 7361 17828 7395
rect 17776 7352 17828 7361
rect 18696 7420 18748 7472
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 9404 7327 9456 7336
rect 9404 7293 9413 7327
rect 9413 7293 9447 7327
rect 9447 7293 9456 7327
rect 9404 7284 9456 7293
rect 9680 7327 9732 7336
rect 9680 7293 9689 7327
rect 9689 7293 9723 7327
rect 9723 7293 9732 7327
rect 9680 7284 9732 7293
rect 11520 7327 11572 7336
rect 11520 7293 11529 7327
rect 11529 7293 11563 7327
rect 11563 7293 11572 7327
rect 11520 7284 11572 7293
rect 14280 7284 14332 7336
rect 15384 7284 15436 7336
rect 13544 7216 13596 7268
rect 18696 7284 18748 7336
rect 19432 7284 19484 7336
rect 20628 7352 20680 7404
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 22928 7463 22980 7472
rect 22928 7429 22937 7463
rect 22937 7429 22971 7463
rect 22971 7429 22980 7463
rect 22928 7420 22980 7429
rect 23112 7488 23164 7540
rect 26424 7488 26476 7540
rect 26608 7531 26660 7540
rect 26608 7497 26617 7531
rect 26617 7497 26651 7531
rect 26651 7497 26660 7531
rect 26608 7488 26660 7497
rect 27528 7488 27580 7540
rect 27620 7488 27672 7540
rect 27712 7488 27764 7540
rect 21088 7284 21140 7336
rect 21272 7284 21324 7336
rect 23572 7352 23624 7404
rect 24032 7395 24084 7404
rect 24032 7361 24041 7395
rect 24041 7361 24075 7395
rect 24075 7361 24084 7395
rect 24032 7352 24084 7361
rect 25044 7420 25096 7472
rect 25320 7420 25372 7472
rect 26240 7420 26292 7472
rect 26332 7420 26384 7472
rect 24492 7395 24544 7404
rect 24492 7361 24501 7395
rect 24501 7361 24535 7395
rect 24535 7361 24544 7395
rect 24492 7352 24544 7361
rect 24584 7352 24636 7404
rect 25228 7352 25280 7404
rect 27344 7420 27396 7472
rect 22008 7216 22060 7268
rect 25412 7284 25464 7336
rect 28540 7352 28592 7404
rect 29000 7395 29052 7404
rect 29000 7361 29009 7395
rect 29009 7361 29043 7395
rect 29043 7361 29052 7395
rect 29000 7352 29052 7361
rect 28264 7327 28316 7336
rect 28264 7293 28273 7327
rect 28273 7293 28307 7327
rect 28307 7293 28316 7327
rect 28264 7284 28316 7293
rect 23572 7216 23624 7268
rect 6184 7148 6236 7200
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11152 7148 11204 7157
rect 12900 7148 12952 7200
rect 13360 7148 13412 7200
rect 14924 7148 14976 7200
rect 15476 7148 15528 7200
rect 15568 7148 15620 7200
rect 17868 7191 17920 7200
rect 17868 7157 17877 7191
rect 17877 7157 17911 7191
rect 17911 7157 17920 7191
rect 17868 7148 17920 7157
rect 18052 7148 18104 7200
rect 20536 7148 20588 7200
rect 20904 7148 20956 7200
rect 24492 7148 24544 7200
rect 24860 7191 24912 7200
rect 24860 7157 24869 7191
rect 24869 7157 24903 7191
rect 24903 7157 24912 7191
rect 24860 7148 24912 7157
rect 25044 7148 25096 7200
rect 25136 7191 25188 7200
rect 25136 7157 25145 7191
rect 25145 7157 25179 7191
rect 25179 7157 25188 7191
rect 25136 7148 25188 7157
rect 26700 7148 26752 7200
rect 27712 7148 27764 7200
rect 28080 7216 28132 7268
rect 29184 7352 29236 7404
rect 29644 7488 29696 7540
rect 30012 7488 30064 7540
rect 31208 7488 31260 7540
rect 31576 7420 31628 7472
rect 30656 7352 30708 7404
rect 31392 7395 31444 7404
rect 31392 7361 31401 7395
rect 31401 7361 31435 7395
rect 31435 7361 31444 7395
rect 31392 7352 31444 7361
rect 31760 7395 31812 7404
rect 31760 7361 31769 7395
rect 31769 7361 31803 7395
rect 31803 7361 31812 7395
rect 31760 7352 31812 7361
rect 31300 7327 31352 7336
rect 31300 7293 31309 7327
rect 31309 7293 31343 7327
rect 31343 7293 31352 7327
rect 31300 7284 31352 7293
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 6000 6987 6052 6996
rect 6000 6953 6009 6987
rect 6009 6953 6043 6987
rect 6043 6953 6052 6987
rect 6000 6944 6052 6953
rect 12348 6987 12400 6996
rect 12348 6953 12357 6987
rect 12357 6953 12391 6987
rect 12391 6953 12400 6987
rect 12348 6944 12400 6953
rect 12808 6987 12860 6996
rect 12808 6953 12817 6987
rect 12817 6953 12851 6987
rect 12851 6953 12860 6987
rect 12808 6944 12860 6953
rect 13636 6944 13688 6996
rect 15568 6944 15620 6996
rect 17776 6944 17828 6996
rect 18052 6987 18104 6996
rect 18052 6953 18061 6987
rect 18061 6953 18095 6987
rect 18095 6953 18104 6987
rect 18052 6944 18104 6953
rect 21272 6944 21324 6996
rect 22468 6944 22520 6996
rect 25412 6987 25464 6996
rect 25412 6953 25421 6987
rect 25421 6953 25455 6987
rect 25455 6953 25464 6987
rect 25412 6944 25464 6953
rect 11152 6876 11204 6928
rect 4620 6808 4672 6860
rect 5080 6808 5132 6860
rect 17316 6876 17368 6928
rect 13728 6808 13780 6860
rect 15752 6808 15804 6860
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 8208 6740 8260 6792
rect 9496 6740 9548 6792
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 15200 6783 15252 6792
rect 15200 6749 15209 6783
rect 15209 6749 15243 6783
rect 15243 6749 15252 6783
rect 15200 6740 15252 6749
rect 4528 6715 4580 6724
rect 4528 6681 4537 6715
rect 4537 6681 4571 6715
rect 4571 6681 4580 6715
rect 4528 6672 4580 6681
rect 6460 6672 6512 6724
rect 16764 6672 16816 6724
rect 18236 6740 18288 6792
rect 19984 6851 20036 6860
rect 19984 6817 19993 6851
rect 19993 6817 20027 6851
rect 20027 6817 20036 6851
rect 19984 6808 20036 6817
rect 24860 6851 24912 6860
rect 24860 6817 24869 6851
rect 24869 6817 24903 6851
rect 24903 6817 24912 6851
rect 24860 6808 24912 6817
rect 18604 6740 18656 6792
rect 18972 6740 19024 6792
rect 20628 6740 20680 6792
rect 21272 6783 21324 6792
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 21364 6740 21416 6792
rect 24952 6783 25004 6792
rect 24952 6749 24961 6783
rect 24961 6749 24995 6783
rect 24995 6749 25004 6783
rect 24952 6740 25004 6749
rect 25596 6783 25648 6792
rect 25596 6749 25605 6783
rect 25605 6749 25639 6783
rect 25639 6749 25648 6783
rect 25596 6740 25648 6749
rect 22100 6672 22152 6724
rect 25412 6715 25464 6724
rect 25412 6681 25421 6715
rect 25421 6681 25455 6715
rect 25455 6681 25464 6715
rect 26056 6740 26108 6792
rect 26240 6783 26292 6792
rect 26240 6749 26249 6783
rect 26249 6749 26283 6783
rect 26283 6749 26292 6783
rect 26240 6740 26292 6749
rect 26608 6944 26660 6996
rect 28724 6944 28776 6996
rect 28908 6944 28960 6996
rect 30932 6944 30984 6996
rect 31300 6944 31352 6996
rect 31392 6944 31444 6996
rect 27896 6876 27948 6928
rect 25412 6672 25464 6681
rect 8484 6604 8536 6656
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 9036 6604 9088 6613
rect 13820 6604 13872 6656
rect 22376 6604 22428 6656
rect 25320 6647 25372 6656
rect 25320 6613 25329 6647
rect 25329 6613 25363 6647
rect 25363 6613 25372 6647
rect 25320 6604 25372 6613
rect 25596 6604 25648 6656
rect 27804 6808 27856 6860
rect 26976 6783 27028 6792
rect 26976 6749 26985 6783
rect 26985 6749 27019 6783
rect 27019 6749 27028 6783
rect 26976 6740 27028 6749
rect 27712 6740 27764 6792
rect 28448 6808 28500 6860
rect 28540 6851 28592 6860
rect 28540 6817 28549 6851
rect 28549 6817 28583 6851
rect 28583 6817 28592 6851
rect 28540 6808 28592 6817
rect 32588 6851 32640 6860
rect 32588 6817 32597 6851
rect 32597 6817 32631 6851
rect 32631 6817 32640 6851
rect 32588 6808 32640 6817
rect 32864 6808 32916 6860
rect 33140 6851 33192 6860
rect 33140 6817 33149 6851
rect 33149 6817 33183 6851
rect 33183 6817 33192 6851
rect 33140 6808 33192 6817
rect 27988 6783 28040 6792
rect 27988 6749 28002 6783
rect 28002 6749 28036 6783
rect 28036 6749 28040 6783
rect 27988 6740 28040 6749
rect 28172 6740 28224 6792
rect 28264 6783 28316 6792
rect 28264 6749 28273 6783
rect 28273 6749 28307 6783
rect 28307 6749 28316 6783
rect 28264 6740 28316 6749
rect 28080 6672 28132 6724
rect 28724 6783 28776 6792
rect 28724 6749 28733 6783
rect 28733 6749 28767 6783
rect 28767 6749 28776 6783
rect 28724 6740 28776 6749
rect 28816 6740 28868 6792
rect 27436 6604 27488 6656
rect 28356 6604 28408 6656
rect 30472 6740 30524 6792
rect 30564 6740 30616 6792
rect 30840 6783 30892 6792
rect 30840 6749 30849 6783
rect 30849 6749 30883 6783
rect 30883 6749 30892 6783
rect 30840 6740 30892 6749
rect 31760 6783 31812 6792
rect 31760 6749 31769 6783
rect 31769 6749 31803 6783
rect 31803 6749 31812 6783
rect 31760 6740 31812 6749
rect 32128 6783 32180 6792
rect 32128 6749 32137 6783
rect 32137 6749 32171 6783
rect 32171 6749 32180 6783
rect 32128 6740 32180 6749
rect 32680 6783 32732 6792
rect 32680 6749 32689 6783
rect 32689 6749 32723 6783
rect 32723 6749 32732 6783
rect 32680 6740 32732 6749
rect 33048 6740 33100 6792
rect 34428 6672 34480 6724
rect 31944 6604 31996 6656
rect 32220 6604 32272 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4528 6400 4580 6452
rect 5172 6400 5224 6452
rect 9496 6400 9548 6452
rect 13912 6400 13964 6452
rect 8852 6332 8904 6384
rect 9404 6332 9456 6384
rect 8208 6264 8260 6316
rect 7472 6196 7524 6248
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 10232 6264 10284 6316
rect 13636 6307 13688 6316
rect 9772 6196 9824 6248
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 14648 6332 14700 6384
rect 17868 6400 17920 6452
rect 18696 6443 18748 6452
rect 18696 6409 18705 6443
rect 18705 6409 18739 6443
rect 18739 6409 18748 6443
rect 18696 6400 18748 6409
rect 19340 6400 19392 6452
rect 19984 6400 20036 6452
rect 20076 6400 20128 6452
rect 23296 6400 23348 6452
rect 12624 6196 12676 6248
rect 12348 6128 12400 6180
rect 7380 6103 7432 6112
rect 7380 6069 7389 6103
rect 7389 6069 7423 6103
rect 7423 6069 7432 6103
rect 7380 6060 7432 6069
rect 8208 6103 8260 6112
rect 8208 6069 8217 6103
rect 8217 6069 8251 6103
rect 8251 6069 8260 6103
rect 8208 6060 8260 6069
rect 8852 6060 8904 6112
rect 9496 6060 9548 6112
rect 15292 6264 15344 6316
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 18144 6264 18196 6316
rect 18604 6332 18656 6384
rect 18972 6264 19024 6316
rect 19708 6307 19760 6316
rect 19708 6273 19717 6307
rect 19717 6273 19751 6307
rect 19751 6273 19760 6307
rect 19708 6264 19760 6273
rect 22560 6332 22612 6384
rect 22928 6332 22980 6384
rect 24952 6400 25004 6452
rect 25228 6400 25280 6452
rect 27988 6443 28040 6452
rect 27988 6409 27997 6443
rect 27997 6409 28031 6443
rect 28031 6409 28040 6443
rect 27988 6400 28040 6409
rect 28172 6443 28224 6452
rect 28172 6409 28181 6443
rect 28181 6409 28215 6443
rect 28215 6409 28224 6443
rect 28172 6400 28224 6409
rect 31024 6400 31076 6452
rect 24492 6332 24544 6384
rect 18144 6171 18196 6180
rect 18144 6137 18153 6171
rect 18153 6137 18187 6171
rect 18187 6137 18196 6171
rect 18144 6128 18196 6137
rect 15200 6060 15252 6112
rect 15384 6060 15436 6112
rect 16488 6060 16540 6112
rect 22652 6264 22704 6316
rect 23112 6264 23164 6316
rect 23572 6307 23624 6316
rect 23572 6273 23581 6307
rect 23581 6273 23615 6307
rect 23615 6273 23624 6307
rect 23572 6264 23624 6273
rect 24032 6264 24084 6316
rect 25320 6332 25372 6384
rect 33140 6400 33192 6452
rect 26056 6264 26108 6316
rect 27804 6307 27856 6316
rect 26792 6196 26844 6248
rect 19524 6060 19576 6112
rect 23020 6103 23072 6112
rect 23020 6069 23029 6103
rect 23029 6069 23063 6103
rect 23063 6069 23072 6103
rect 23020 6060 23072 6069
rect 24400 6128 24452 6180
rect 27804 6273 27813 6307
rect 27813 6273 27847 6307
rect 27847 6273 27856 6307
rect 27804 6264 27856 6273
rect 27620 6196 27672 6248
rect 27436 6128 27488 6180
rect 32220 6264 32272 6316
rect 32680 6264 32732 6316
rect 32588 6128 32640 6180
rect 32772 6171 32824 6180
rect 32772 6137 32781 6171
rect 32781 6137 32815 6171
rect 32815 6137 32824 6171
rect 32772 6128 32824 6137
rect 27620 6103 27672 6112
rect 27620 6069 27629 6103
rect 27629 6069 27663 6103
rect 27663 6069 27672 6103
rect 27620 6060 27672 6069
rect 27804 6060 27856 6112
rect 28908 6060 28960 6112
rect 32036 6060 32088 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 8208 5856 8260 5908
rect 5080 5763 5132 5772
rect 5080 5729 5089 5763
rect 5089 5729 5123 5763
rect 5123 5729 5132 5763
rect 6920 5763 6972 5772
rect 5080 5720 5132 5729
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 9312 5856 9364 5908
rect 10324 5856 10376 5908
rect 14188 5856 14240 5908
rect 15476 5856 15528 5908
rect 16304 5856 16356 5908
rect 18144 5856 18196 5908
rect 9680 5788 9732 5840
rect 6460 5652 6512 5704
rect 8484 5652 8536 5704
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 9496 5695 9548 5704
rect 9496 5661 9506 5695
rect 9506 5661 9540 5695
rect 9540 5661 9548 5695
rect 9496 5652 9548 5661
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 10324 5695 10376 5704
rect 10324 5661 10331 5695
rect 10331 5661 10376 5695
rect 5632 5584 5684 5636
rect 10324 5652 10376 5661
rect 13544 5788 13596 5840
rect 14924 5763 14976 5772
rect 12440 5652 12492 5704
rect 8208 5516 8260 5568
rect 10416 5627 10468 5636
rect 10416 5593 10425 5627
rect 10425 5593 10459 5627
rect 10459 5593 10468 5627
rect 10416 5584 10468 5593
rect 12624 5652 12676 5704
rect 14924 5729 14933 5763
rect 14933 5729 14967 5763
rect 14967 5729 14976 5763
rect 14924 5720 14976 5729
rect 12992 5584 13044 5636
rect 15200 5652 15252 5704
rect 15752 5720 15804 5772
rect 17132 5695 17184 5704
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 20076 5856 20128 5908
rect 22836 5856 22888 5908
rect 23204 5856 23256 5908
rect 27436 5856 27488 5908
rect 30472 5899 30524 5908
rect 30472 5865 30481 5899
rect 30481 5865 30515 5899
rect 30515 5865 30524 5899
rect 30472 5856 30524 5865
rect 32036 5899 32088 5908
rect 32036 5865 32045 5899
rect 32045 5865 32079 5899
rect 32079 5865 32088 5899
rect 32036 5856 32088 5865
rect 32220 5899 32272 5908
rect 32220 5865 32229 5899
rect 32229 5865 32263 5899
rect 32263 5865 32272 5899
rect 32220 5856 32272 5865
rect 24676 5788 24728 5840
rect 19340 5720 19392 5772
rect 19524 5720 19576 5772
rect 20076 5695 20128 5704
rect 20076 5661 20085 5695
rect 20085 5661 20119 5695
rect 20119 5661 20128 5695
rect 20076 5652 20128 5661
rect 20444 5695 20496 5704
rect 20444 5661 20453 5695
rect 20453 5661 20487 5695
rect 20487 5661 20496 5695
rect 20444 5652 20496 5661
rect 20536 5652 20588 5704
rect 14280 5584 14332 5636
rect 15936 5584 15988 5636
rect 16120 5584 16172 5636
rect 19708 5584 19760 5636
rect 22652 5652 22704 5704
rect 22928 5695 22980 5704
rect 22928 5661 22937 5695
rect 22937 5661 22971 5695
rect 22971 5661 22980 5695
rect 22928 5652 22980 5661
rect 23112 5695 23164 5704
rect 23112 5661 23121 5695
rect 23121 5661 23155 5695
rect 23155 5661 23164 5695
rect 23112 5652 23164 5661
rect 23572 5695 23624 5704
rect 23572 5661 23581 5695
rect 23581 5661 23615 5695
rect 23615 5661 23624 5695
rect 23572 5652 23624 5661
rect 23664 5695 23716 5704
rect 23664 5661 23673 5695
rect 23673 5661 23707 5695
rect 23707 5661 23716 5695
rect 23664 5652 23716 5661
rect 24400 5652 24452 5704
rect 24952 5720 25004 5772
rect 28356 5788 28408 5840
rect 29276 5788 29328 5840
rect 29184 5720 29236 5772
rect 31760 5652 31812 5704
rect 32128 5695 32180 5704
rect 32128 5661 32137 5695
rect 32137 5661 32171 5695
rect 32171 5661 32180 5695
rect 32128 5652 32180 5661
rect 9864 5516 9916 5568
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 11704 5516 11756 5568
rect 13636 5516 13688 5568
rect 13820 5559 13872 5568
rect 13820 5525 13829 5559
rect 13829 5525 13863 5559
rect 13863 5525 13872 5559
rect 13820 5516 13872 5525
rect 14372 5559 14424 5568
rect 14372 5525 14381 5559
rect 14381 5525 14415 5559
rect 14415 5525 14424 5559
rect 14372 5516 14424 5525
rect 15384 5516 15436 5568
rect 19984 5516 20036 5568
rect 20996 5516 21048 5568
rect 22836 5516 22888 5568
rect 30196 5584 30248 5636
rect 30288 5627 30340 5636
rect 30288 5593 30297 5627
rect 30297 5593 30331 5627
rect 30331 5593 30340 5627
rect 30288 5584 30340 5593
rect 24400 5559 24452 5568
rect 24400 5525 24409 5559
rect 24409 5525 24443 5559
rect 24443 5525 24452 5559
rect 24400 5516 24452 5525
rect 29828 5516 29880 5568
rect 31944 5584 31996 5636
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 5632 5312 5684 5364
rect 7380 5312 7432 5364
rect 8852 5355 8904 5364
rect 8852 5321 8861 5355
rect 8861 5321 8895 5355
rect 8895 5321 8904 5355
rect 8852 5312 8904 5321
rect 8208 5219 8260 5228
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 8208 5176 8260 5185
rect 9036 5176 9088 5228
rect 9864 5312 9916 5364
rect 11520 5312 11572 5364
rect 12164 5312 12216 5364
rect 9864 5176 9916 5228
rect 10416 5244 10468 5296
rect 10048 5176 10100 5228
rect 11704 5244 11756 5296
rect 12532 5244 12584 5296
rect 15200 5355 15252 5364
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 17132 5312 17184 5364
rect 20168 5312 20220 5364
rect 20444 5312 20496 5364
rect 22836 5312 22888 5364
rect 23572 5312 23624 5364
rect 23664 5355 23716 5364
rect 23664 5321 23673 5355
rect 23673 5321 23707 5355
rect 23707 5321 23716 5355
rect 23664 5312 23716 5321
rect 24860 5312 24912 5364
rect 13636 5244 13688 5296
rect 19340 5287 19392 5296
rect 19340 5253 19349 5287
rect 19349 5253 19383 5287
rect 19383 5253 19392 5287
rect 19340 5244 19392 5253
rect 19432 5244 19484 5296
rect 9680 5108 9732 5160
rect 12992 5108 13044 5160
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 12532 4972 12584 5024
rect 16120 5176 16172 5228
rect 20996 5244 21048 5296
rect 20904 5219 20956 5228
rect 20904 5185 20913 5219
rect 20913 5185 20947 5219
rect 20947 5185 20956 5219
rect 20904 5176 20956 5185
rect 22744 5176 22796 5228
rect 23020 5219 23072 5228
rect 23020 5185 23029 5219
rect 23029 5185 23063 5219
rect 23063 5185 23072 5219
rect 23020 5176 23072 5185
rect 23112 5176 23164 5228
rect 23204 5219 23256 5228
rect 23204 5185 23213 5219
rect 23213 5185 23247 5219
rect 23247 5185 23256 5219
rect 23204 5176 23256 5185
rect 15384 5108 15436 5160
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 16672 5151 16724 5160
rect 16672 5117 16681 5151
rect 16681 5117 16715 5151
rect 16715 5117 16724 5151
rect 16672 5108 16724 5117
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 22376 5108 22428 5117
rect 23296 5040 23348 5092
rect 24676 5176 24728 5228
rect 25412 5176 25464 5228
rect 27620 5312 27672 5364
rect 26240 5176 26292 5228
rect 28448 5244 28500 5296
rect 27620 5219 27672 5228
rect 27620 5185 27629 5219
rect 27629 5185 27663 5219
rect 27663 5185 27672 5219
rect 27620 5176 27672 5185
rect 27712 5219 27764 5228
rect 27712 5185 27721 5219
rect 27721 5185 27755 5219
rect 27755 5185 27764 5219
rect 27712 5176 27764 5185
rect 24400 5108 24452 5160
rect 26976 5108 27028 5160
rect 29276 5176 29328 5228
rect 28264 5108 28316 5160
rect 26056 5040 26108 5092
rect 29184 5040 29236 5092
rect 16396 5015 16448 5024
rect 16396 4981 16405 5015
rect 16405 4981 16439 5015
rect 16439 4981 16448 5015
rect 16396 4972 16448 4981
rect 23388 4972 23440 5024
rect 24400 4972 24452 5024
rect 29644 4972 29696 5024
rect 29828 5176 29880 5228
rect 30288 5312 30340 5364
rect 32128 5312 32180 5364
rect 30104 5176 30156 5228
rect 29828 5083 29880 5092
rect 29828 5049 29837 5083
rect 29837 5049 29871 5083
rect 29871 5049 29880 5083
rect 29828 5040 29880 5049
rect 30012 4972 30064 5024
rect 30288 5015 30340 5024
rect 30288 4981 30297 5015
rect 30297 4981 30331 5015
rect 30331 4981 30340 5015
rect 30288 4972 30340 4981
rect 30656 5083 30708 5092
rect 30656 5049 30665 5083
rect 30665 5049 30699 5083
rect 30699 5049 30708 5083
rect 30656 5040 30708 5049
rect 31760 5176 31812 5228
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 11152 4768 11204 4820
rect 12624 4768 12676 4820
rect 15844 4768 15896 4820
rect 16396 4768 16448 4820
rect 16672 4768 16724 4820
rect 19984 4768 20036 4820
rect 20168 4811 20220 4820
rect 20168 4777 20177 4811
rect 20177 4777 20211 4811
rect 20211 4777 20220 4811
rect 20168 4768 20220 4777
rect 20904 4768 20956 4820
rect 20996 4768 21048 4820
rect 12164 4632 12216 4684
rect 23388 4768 23440 4820
rect 24400 4811 24452 4820
rect 24400 4777 24409 4811
rect 24409 4777 24443 4811
rect 24443 4777 24452 4811
rect 24400 4768 24452 4777
rect 25504 4768 25556 4820
rect 26056 4811 26108 4820
rect 26056 4777 26065 4811
rect 26065 4777 26099 4811
rect 26099 4777 26108 4811
rect 26056 4768 26108 4777
rect 27620 4768 27672 4820
rect 29184 4768 29236 4820
rect 30012 4811 30064 4820
rect 30012 4777 30021 4811
rect 30021 4777 30055 4811
rect 30055 4777 30064 4811
rect 30012 4768 30064 4777
rect 30196 4768 30248 4820
rect 3884 4564 3936 4616
rect 9772 4564 9824 4616
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 15936 4564 15988 4616
rect 20260 4632 20312 4684
rect 27896 4700 27948 4752
rect 29828 4700 29880 4752
rect 30656 4700 30708 4752
rect 16304 4607 16356 4616
rect 16304 4573 16313 4607
rect 16313 4573 16347 4607
rect 16347 4573 16356 4607
rect 16304 4564 16356 4573
rect 16488 4564 16540 4616
rect 20352 4564 20404 4616
rect 21824 4607 21876 4616
rect 21824 4573 21833 4607
rect 21833 4573 21867 4607
rect 21867 4573 21876 4607
rect 21824 4564 21876 4573
rect 23480 4632 23532 4684
rect 940 4496 992 4548
rect 12532 4496 12584 4548
rect 14464 4539 14516 4548
rect 14464 4505 14473 4539
rect 14473 4505 14507 4539
rect 14507 4505 14516 4539
rect 14464 4496 14516 4505
rect 16764 4428 16816 4480
rect 20076 4496 20128 4548
rect 20536 4496 20588 4548
rect 22744 4496 22796 4548
rect 23296 4539 23348 4548
rect 23296 4505 23305 4539
rect 23305 4505 23339 4539
rect 23339 4505 23348 4539
rect 23296 4496 23348 4505
rect 24492 4496 24544 4548
rect 24860 4607 24912 4616
rect 24860 4573 24869 4607
rect 24869 4573 24903 4607
rect 24903 4573 24912 4607
rect 24860 4564 24912 4573
rect 25412 4632 25464 4684
rect 24676 4496 24728 4548
rect 25596 4607 25648 4616
rect 25596 4573 25605 4607
rect 25605 4573 25639 4607
rect 25639 4573 25648 4607
rect 25596 4564 25648 4573
rect 26976 4632 27028 4684
rect 26332 4607 26384 4616
rect 26332 4573 26341 4607
rect 26341 4573 26375 4607
rect 26375 4573 26384 4607
rect 27988 4675 28040 4684
rect 27988 4641 27997 4675
rect 27997 4641 28031 4675
rect 28031 4641 28040 4675
rect 27988 4632 28040 4641
rect 28080 4632 28132 4684
rect 29276 4632 29328 4684
rect 26332 4564 26384 4573
rect 29644 4564 29696 4616
rect 30288 4607 30340 4616
rect 30288 4573 30297 4607
rect 30297 4573 30331 4607
rect 30331 4573 30340 4607
rect 30288 4564 30340 4573
rect 31760 4496 31812 4548
rect 27712 4428 27764 4480
rect 31944 4428 31996 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 9128 4224 9180 4276
rect 9680 4224 9732 4276
rect 14464 4224 14516 4276
rect 25504 4224 25556 4276
rect 27988 4224 28040 4276
rect 8576 4156 8628 4208
rect 6920 4088 6972 4140
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 25136 4131 25188 4140
rect 25136 4097 25145 4131
rect 25145 4097 25179 4131
rect 25179 4097 25188 4131
rect 25136 4088 25188 4097
rect 25228 4131 25280 4140
rect 25228 4097 25237 4131
rect 25237 4097 25271 4131
rect 25271 4097 25280 4131
rect 25228 4088 25280 4097
rect 26332 4020 26384 4072
rect 27896 4088 27948 4140
rect 30104 4088 30156 4140
rect 25412 3952 25464 4004
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 17224 3136 17276 3188
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 12532 3043 12584 3052
rect 12532 3009 12541 3043
rect 12541 3009 12575 3043
rect 12575 3009 12584 3043
rect 12532 3000 12584 3009
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 15108 3043 15160 3052
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 37556 3111 37608 3120
rect 37556 3077 37565 3111
rect 37565 3077 37599 3111
rect 37599 3077 37608 3111
rect 37556 3068 37608 3077
rect 25964 3000 26016 3052
rect 1768 2839 1820 2848
rect 1768 2805 1777 2839
rect 1777 2805 1811 2839
rect 1811 2805 1820 2839
rect 1768 2796 1820 2805
rect 2228 2839 2280 2848
rect 2228 2805 2237 2839
rect 2237 2805 2271 2839
rect 2271 2805 2280 2839
rect 2228 2796 2280 2805
rect 8392 2796 8444 2848
rect 12992 2839 13044 2848
rect 12992 2805 13001 2839
rect 13001 2805 13035 2839
rect 13035 2805 13044 2839
rect 12992 2796 13044 2805
rect 14924 2839 14976 2848
rect 14924 2805 14933 2839
rect 14933 2805 14967 2839
rect 14967 2805 14976 2839
rect 14924 2796 14976 2805
rect 17408 2839 17460 2848
rect 17408 2805 17417 2839
rect 17417 2805 17451 2839
rect 17451 2805 17460 2839
rect 17408 2796 17460 2805
rect 19800 2839 19852 2848
rect 19800 2805 19809 2839
rect 19809 2805 19843 2839
rect 19843 2805 19852 2839
rect 19800 2796 19852 2805
rect 37188 2796 37240 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 8760 2592 8812 2644
rect 10140 2592 10192 2644
rect 8944 2456 8996 2508
rect 1768 2431 1820 2440
rect 1768 2397 1777 2431
rect 1777 2397 1811 2431
rect 1811 2397 1820 2431
rect 1768 2388 1820 2397
rect 2228 2388 2280 2440
rect 4804 2388 4856 2440
rect 8392 2388 8444 2440
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 12992 2388 13044 2440
rect 14924 2388 14976 2440
rect 17408 2388 17460 2440
rect 19800 2431 19852 2440
rect 19800 2397 19809 2431
rect 19809 2397 19843 2431
rect 19843 2397 19852 2431
rect 19800 2388 19852 2397
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 20 2320 72 2372
rect 2044 2363 2096 2372
rect 2044 2329 2053 2363
rect 2053 2329 2087 2363
rect 2087 2329 2096 2363
rect 2044 2320 2096 2329
rect 3976 2363 4028 2372
rect 3976 2329 3985 2363
rect 3985 2329 4019 2363
rect 4019 2329 4028 2363
rect 3976 2320 4028 2329
rect 6552 2363 6604 2372
rect 6552 2329 6561 2363
rect 6561 2329 6595 2363
rect 6595 2329 6604 2363
rect 6552 2320 6604 2329
rect 10968 2320 11020 2372
rect 14648 2320 14700 2372
rect 12900 2252 12952 2304
rect 15016 2252 15068 2304
rect 17408 2252 17460 2304
rect 19432 2363 19484 2372
rect 19432 2329 19441 2363
rect 19441 2329 19475 2363
rect 19475 2329 19484 2363
rect 19432 2320 19484 2329
rect 26424 2252 26476 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 18 40762 74 41562
rect 1950 40762 2006 41562
rect 4526 40882 4582 41562
rect 4526 40854 4936 40882
rect 4526 40762 4582 40854
rect 32 39098 60 40762
rect 4908 39098 4936 40854
rect 6458 40762 6514 41562
rect 9034 40762 9090 41562
rect 10966 40762 11022 41562
rect 12898 40882 12954 41562
rect 12898 40854 13216 40882
rect 12898 40762 12954 40854
rect 9048 39098 9076 40762
rect 10980 39114 11008 40762
rect 10980 39098 11100 39114
rect 13188 39098 13216 40854
rect 15474 40762 15530 41562
rect 17406 40762 17462 41562
rect 19982 40882 20038 41562
rect 19982 40854 20116 40882
rect 19982 40762 20038 40854
rect 20 39092 72 39098
rect 20 39034 72 39040
rect 4896 39092 4948 39098
rect 4896 39034 4948 39040
rect 9036 39092 9088 39098
rect 10980 39092 11112 39098
rect 10980 39086 11060 39092
rect 9036 39034 9088 39040
rect 11060 39034 11112 39040
rect 13176 39092 13228 39098
rect 13176 39034 13228 39040
rect 15488 39030 15516 40762
rect 17420 39098 17448 40762
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 17408 39092 17460 39098
rect 17408 39034 17460 39040
rect 12348 39024 12400 39030
rect 12348 38966 12400 38972
rect 15476 39024 15528 39030
rect 15476 38966 15528 38972
rect 1768 38956 1820 38962
rect 1768 38898 1820 38904
rect 5080 38956 5132 38962
rect 5080 38898 5132 38904
rect 9220 38956 9272 38962
rect 9220 38898 9272 38904
rect 12072 38956 12124 38962
rect 12072 38898 12124 38904
rect 940 37188 992 37194
rect 940 37130 992 37136
rect 952 36825 980 37130
rect 938 36816 994 36825
rect 938 36751 994 36760
rect 1780 35894 1808 38898
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 5092 38554 5120 38898
rect 9232 38554 9260 38898
rect 5080 38548 5132 38554
rect 5080 38490 5132 38496
rect 9220 38548 9272 38554
rect 9220 38490 9272 38496
rect 5170 38448 5226 38457
rect 5170 38383 5226 38392
rect 5184 38350 5212 38383
rect 5172 38344 5224 38350
rect 5172 38286 5224 38292
rect 8576 38344 8628 38350
rect 8576 38286 8628 38292
rect 9036 38344 9088 38350
rect 9036 38286 9088 38292
rect 11336 38344 11388 38350
rect 11336 38286 11388 38292
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 8300 37256 8352 37262
rect 8300 37198 8352 37204
rect 7196 37188 7248 37194
rect 7196 37130 7248 37136
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 6828 36236 6880 36242
rect 6828 36178 6880 36184
rect 5724 36168 5776 36174
rect 5724 36110 5776 36116
rect 1780 35866 2176 35894
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 940 25696 992 25702
rect 940 25638 992 25644
rect 952 25265 980 25638
rect 1400 25288 1452 25294
rect 938 25256 994 25265
rect 1400 25230 1452 25236
rect 938 25191 994 25200
rect 1412 24750 1440 25230
rect 1400 24744 1452 24750
rect 1400 24686 1452 24692
rect 1676 24744 1728 24750
rect 1676 24686 1728 24692
rect 1412 24342 1440 24686
rect 1688 24410 1716 24686
rect 1676 24404 1728 24410
rect 1676 24346 1728 24352
rect 1400 24336 1452 24342
rect 1400 24278 1452 24284
rect 1412 21486 1440 24278
rect 1780 23322 1808 25842
rect 1860 25832 1912 25838
rect 1860 25774 1912 25780
rect 1872 25294 1900 25774
rect 1860 25288 1912 25294
rect 1860 25230 1912 25236
rect 1952 23860 2004 23866
rect 1952 23802 2004 23808
rect 1768 23316 1820 23322
rect 1768 23258 1820 23264
rect 1964 23118 1992 23802
rect 1952 23112 2004 23118
rect 1952 23054 2004 23060
rect 1860 22976 1912 22982
rect 1860 22918 1912 22924
rect 1768 21888 1820 21894
rect 1768 21830 1820 21836
rect 1780 21690 1808 21830
rect 1768 21684 1820 21690
rect 1768 21626 1820 21632
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 19514 1440 21422
rect 1872 20942 1900 22918
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 1964 21690 1992 21966
rect 1952 21684 2004 21690
rect 1952 21626 2004 21632
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1504 20641 1532 20742
rect 1490 20632 1546 20641
rect 1490 20567 1546 20576
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 1400 19508 1452 19514
rect 1400 19450 1452 19456
rect 1780 19446 1808 19654
rect 1768 19440 1820 19446
rect 1768 19382 1820 19388
rect 940 18692 992 18698
rect 940 18634 992 18640
rect 1768 18692 1820 18698
rect 1768 18634 1820 18640
rect 952 18465 980 18634
rect 938 18456 994 18465
rect 938 18391 994 18400
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1688 17746 1716 18158
rect 1780 17882 1808 18634
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1964 17678 1992 18566
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 2056 17678 2084 18022
rect 2148 17882 2176 35866
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 5540 34604 5592 34610
rect 5540 34546 5592 34552
rect 5356 34400 5408 34406
rect 5356 34342 5408 34348
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 5368 33930 5396 34342
rect 5356 33924 5408 33930
rect 5356 33866 5408 33872
rect 5552 33658 5580 34546
rect 5736 34066 5764 36110
rect 6276 36100 6328 36106
rect 6276 36042 6328 36048
rect 6288 35834 6316 36042
rect 6276 35828 6328 35834
rect 6276 35770 6328 35776
rect 5724 34060 5776 34066
rect 5644 34020 5724 34048
rect 5540 33652 5592 33658
rect 5540 33594 5592 33600
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 3976 32904 4028 32910
rect 3976 32846 4028 32852
rect 3988 31822 4016 32846
rect 4896 32836 4948 32842
rect 4896 32778 4948 32784
rect 4908 32570 4936 32778
rect 4896 32564 4948 32570
rect 4896 32506 4948 32512
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3976 31816 4028 31822
rect 3976 31758 4028 31764
rect 3988 30734 4016 31758
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 5644 30734 5672 34020
rect 5724 34002 5776 34008
rect 6840 33998 6868 36178
rect 7208 35170 7236 37130
rect 8312 36922 8340 37198
rect 8300 36916 8352 36922
rect 8300 36858 8352 36864
rect 7472 36576 7524 36582
rect 7472 36518 7524 36524
rect 7484 36242 7512 36518
rect 7472 36236 7524 36242
rect 7472 36178 7524 36184
rect 7748 36032 7800 36038
rect 7748 35974 7800 35980
rect 7760 35834 7788 35974
rect 7748 35828 7800 35834
rect 7748 35770 7800 35776
rect 8116 35828 8168 35834
rect 8116 35770 8168 35776
rect 7472 35624 7524 35630
rect 7472 35566 7524 35572
rect 7208 35154 7328 35170
rect 7196 35148 7328 35154
rect 7248 35142 7328 35148
rect 7196 35090 7248 35096
rect 7196 35012 7248 35018
rect 7196 34954 7248 34960
rect 7208 34746 7236 34954
rect 7196 34740 7248 34746
rect 7196 34682 7248 34688
rect 7300 33998 7328 35142
rect 6368 33992 6420 33998
rect 6368 33934 6420 33940
rect 6828 33992 6880 33998
rect 6828 33934 6880 33940
rect 7288 33992 7340 33998
rect 7288 33934 7340 33940
rect 5908 33448 5960 33454
rect 5908 33390 5960 33396
rect 5920 32910 5948 33390
rect 6380 33046 6408 33934
rect 6736 33856 6788 33862
rect 6736 33798 6788 33804
rect 7196 33856 7248 33862
rect 7196 33798 7248 33804
rect 6748 33658 6776 33798
rect 7208 33658 7236 33798
rect 6736 33652 6788 33658
rect 6736 33594 6788 33600
rect 7196 33652 7248 33658
rect 7196 33594 7248 33600
rect 7300 33538 7328 33934
rect 7208 33510 7328 33538
rect 7208 33114 7236 33510
rect 7288 33448 7340 33454
rect 7288 33390 7340 33396
rect 7300 33114 7328 33390
rect 7484 33318 7512 35566
rect 8128 34678 8156 35770
rect 8208 35624 8260 35630
rect 8208 35566 8260 35572
rect 8300 35624 8352 35630
rect 8300 35566 8352 35572
rect 8220 35086 8248 35566
rect 8312 35086 8340 35566
rect 8208 35080 8260 35086
rect 8208 35022 8260 35028
rect 8300 35080 8352 35086
rect 8300 35022 8352 35028
rect 8116 34672 8168 34678
rect 8116 34614 8168 34620
rect 8220 34610 8248 35022
rect 8208 34604 8260 34610
rect 8208 34546 8260 34552
rect 7472 33312 7524 33318
rect 7472 33254 7524 33260
rect 7196 33108 7248 33114
rect 7196 33050 7248 33056
rect 7288 33108 7340 33114
rect 7288 33050 7340 33056
rect 6368 33040 6420 33046
rect 6368 32982 6420 32988
rect 5908 32904 5960 32910
rect 5908 32846 5960 32852
rect 6276 32768 6328 32774
rect 6276 32710 6328 32716
rect 6288 32570 6316 32710
rect 6276 32564 6328 32570
rect 6276 32506 6328 32512
rect 5724 32360 5776 32366
rect 5724 32302 5776 32308
rect 5736 31890 5764 32302
rect 5724 31884 5776 31890
rect 5724 31826 5776 31832
rect 3976 30728 4028 30734
rect 3976 30670 4028 30676
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 3988 29646 4016 30670
rect 4252 30592 4304 30598
rect 4252 30534 4304 30540
rect 4264 30190 4292 30534
rect 5264 30320 5316 30326
rect 5264 30262 5316 30268
rect 4252 30184 4304 30190
rect 4252 30126 4304 30132
rect 5276 30054 5304 30262
rect 5264 30048 5316 30054
rect 5264 29990 5316 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3976 29640 4028 29646
rect 3976 29582 4028 29588
rect 4068 29504 4120 29510
rect 4068 29446 4120 29452
rect 4080 29306 4108 29446
rect 4068 29300 4120 29306
rect 4068 29242 4120 29248
rect 5276 29170 5304 29990
rect 5448 29504 5500 29510
rect 5448 29446 5500 29452
rect 5264 29164 5316 29170
rect 5264 29106 5316 29112
rect 4620 28960 4672 28966
rect 4620 28902 4672 28908
rect 5356 28960 5408 28966
rect 5356 28902 5408 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4632 28762 4660 28902
rect 4620 28756 4672 28762
rect 4620 28698 4672 28704
rect 4252 28416 4304 28422
rect 4252 28358 4304 28364
rect 4264 28218 4292 28358
rect 4252 28212 4304 28218
rect 4252 28154 4304 28160
rect 4620 28144 4672 28150
rect 4620 28086 4672 28092
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27674 4660 28086
rect 5368 28082 5396 28902
rect 5460 28558 5488 29446
rect 5644 28558 5672 30670
rect 5736 30054 5764 31826
rect 6380 30938 6408 32982
rect 6828 32972 6880 32978
rect 6828 32914 6880 32920
rect 6552 32904 6604 32910
rect 6552 32846 6604 32852
rect 6564 31822 6592 32846
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6368 30932 6420 30938
rect 6368 30874 6420 30880
rect 6184 30660 6236 30666
rect 6184 30602 6236 30608
rect 6196 30394 6224 30602
rect 6184 30388 6236 30394
rect 6184 30330 6236 30336
rect 6840 30054 6868 32914
rect 7380 32768 7432 32774
rect 7380 32710 7432 32716
rect 7392 31822 7420 32710
rect 7380 31816 7432 31822
rect 7300 31776 7380 31804
rect 7300 30258 7328 31776
rect 7380 31758 7432 31764
rect 7484 30802 7512 33254
rect 8220 32910 8248 34546
rect 8312 33522 8340 35022
rect 8300 33516 8352 33522
rect 8300 33458 8352 33464
rect 7840 32904 7892 32910
rect 7840 32846 7892 32852
rect 8208 32904 8260 32910
rect 8208 32846 8260 32852
rect 7852 32026 7880 32846
rect 8116 32836 8168 32842
rect 8116 32778 8168 32784
rect 8128 32570 8156 32778
rect 8116 32564 8168 32570
rect 8116 32506 8168 32512
rect 7840 32020 7892 32026
rect 7840 31962 7892 31968
rect 7656 31816 7708 31822
rect 8116 31816 8168 31822
rect 7708 31776 7972 31804
rect 7656 31758 7708 31764
rect 7840 31680 7892 31686
rect 7840 31622 7892 31628
rect 7852 31278 7880 31622
rect 7840 31272 7892 31278
rect 7840 31214 7892 31220
rect 7472 30796 7524 30802
rect 7472 30738 7524 30744
rect 7288 30252 7340 30258
rect 7116 30212 7288 30240
rect 5724 30048 5776 30054
rect 5724 29990 5776 29996
rect 6828 30048 6880 30054
rect 6828 29990 6880 29996
rect 6840 29714 6868 29990
rect 6920 29776 6972 29782
rect 6920 29718 6972 29724
rect 6828 29708 6880 29714
rect 6828 29650 6880 29656
rect 6092 29572 6144 29578
rect 6092 29514 6144 29520
rect 6104 29238 6132 29514
rect 6828 29504 6880 29510
rect 6828 29446 6880 29452
rect 6840 29306 6868 29446
rect 6828 29300 6880 29306
rect 6828 29242 6880 29248
rect 6092 29232 6144 29238
rect 6092 29174 6144 29180
rect 6552 28960 6604 28966
rect 6552 28902 6604 28908
rect 6564 28626 6592 28902
rect 6552 28620 6604 28626
rect 6552 28562 6604 28568
rect 5448 28552 5500 28558
rect 5448 28494 5500 28500
rect 5632 28552 5684 28558
rect 5632 28494 5684 28500
rect 6840 28218 6868 29242
rect 6932 29034 6960 29718
rect 7012 29096 7064 29102
rect 7116 29084 7144 30212
rect 7288 30194 7340 30200
rect 7064 29056 7144 29084
rect 7012 29038 7064 29044
rect 6920 29028 6972 29034
rect 6920 28970 6972 28976
rect 6828 28212 6880 28218
rect 6828 28154 6880 28160
rect 5356 28076 5408 28082
rect 5356 28018 5408 28024
rect 6000 28076 6052 28082
rect 6000 28018 6052 28024
rect 4620 27668 4672 27674
rect 4620 27610 4672 27616
rect 4066 27296 4122 27305
rect 4066 27231 4122 27240
rect 3884 26240 3936 26246
rect 3884 26182 3936 26188
rect 3896 25974 3924 26182
rect 3884 25968 3936 25974
rect 3884 25910 3936 25916
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 3056 25900 3108 25906
rect 3056 25842 3108 25848
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 2884 25362 2912 25638
rect 2872 25356 2924 25362
rect 2872 25298 2924 25304
rect 2872 25220 2924 25226
rect 2976 25208 3004 25842
rect 2924 25180 3004 25208
rect 2872 25162 2924 25168
rect 2884 24750 2912 25162
rect 2872 24744 2924 24750
rect 2872 24686 2924 24692
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2792 23322 2820 24006
rect 2780 23316 2832 23322
rect 2780 23258 2832 23264
rect 2884 23202 2912 24686
rect 3068 24410 3096 25842
rect 3608 25832 3660 25838
rect 3608 25774 3660 25780
rect 3620 25498 3648 25774
rect 3608 25492 3660 25498
rect 3608 25434 3660 25440
rect 3148 24608 3200 24614
rect 3148 24550 3200 24556
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3056 24404 3108 24410
rect 3056 24346 3108 24352
rect 3160 24138 3188 24550
rect 3988 24274 4016 24550
rect 4080 24410 4108 27231
rect 6012 26790 6040 28018
rect 6368 27872 6420 27878
rect 6368 27814 6420 27820
rect 6380 27470 6408 27814
rect 6932 27470 6960 28970
rect 6368 27464 6420 27470
rect 6368 27406 6420 27412
rect 6920 27464 6972 27470
rect 6920 27406 6972 27412
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6840 27130 6868 27270
rect 6828 27124 6880 27130
rect 6828 27066 6880 27072
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 5080 26308 5132 26314
rect 5080 26250 5132 26256
rect 5092 26042 5120 26250
rect 6012 26246 6040 26726
rect 6932 26586 6960 26862
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 6000 26240 6052 26246
rect 6000 26182 6052 26188
rect 6920 26240 6972 26246
rect 6920 26182 6972 26188
rect 5080 26036 5132 26042
rect 5080 25978 5132 25984
rect 5080 25696 5132 25702
rect 5080 25638 5132 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4356 24954 4384 25230
rect 4620 25152 4672 25158
rect 4620 25094 4672 25100
rect 4344 24948 4396 24954
rect 4344 24890 4396 24896
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 24404 4120 24410
rect 4068 24346 4120 24352
rect 3240 24268 3292 24274
rect 3240 24210 3292 24216
rect 3976 24268 4028 24274
rect 3976 24210 4028 24216
rect 3148 24132 3200 24138
rect 3148 24074 3200 24080
rect 3160 23202 3188 24074
rect 2792 23174 2912 23202
rect 3068 23174 3188 23202
rect 2688 23112 2740 23118
rect 2688 23054 2740 23060
rect 2504 22976 2556 22982
rect 2504 22918 2556 22924
rect 2516 22710 2544 22918
rect 2700 22778 2728 23054
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2504 22704 2556 22710
rect 2504 22646 2556 22652
rect 2792 21554 2820 23174
rect 2872 22976 2924 22982
rect 2872 22918 2924 22924
rect 2884 22574 2912 22918
rect 3068 22710 3096 23174
rect 3148 23112 3200 23118
rect 3148 23054 3200 23060
rect 3160 22778 3188 23054
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 3056 22704 3108 22710
rect 2962 22672 3018 22681
rect 3056 22646 3108 22652
rect 2962 22607 2964 22616
rect 3016 22607 3018 22616
rect 2964 22578 3016 22584
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2884 20806 2912 22510
rect 3252 22094 3280 24210
rect 3988 23662 4016 24210
rect 4632 24206 4660 25094
rect 5092 24954 5120 25638
rect 5080 24948 5132 24954
rect 5080 24890 5132 24896
rect 5816 24948 5868 24954
rect 5816 24890 5868 24896
rect 4804 24744 4856 24750
rect 4804 24686 4856 24692
rect 4620 24200 4672 24206
rect 4672 24160 4752 24188
rect 4620 24142 4672 24148
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23322 4660 24006
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 4620 23316 4672 23322
rect 4620 23258 4672 23264
rect 3608 23112 3660 23118
rect 3608 23054 3660 23060
rect 3620 22506 3648 23054
rect 3976 22976 4028 22982
rect 3976 22918 4028 22924
rect 3988 22778 4016 22918
rect 3976 22772 4028 22778
rect 3976 22714 4028 22720
rect 3884 22636 3936 22642
rect 3884 22578 3936 22584
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 3608 22500 3660 22506
rect 3608 22442 3660 22448
rect 3700 22432 3752 22438
rect 3700 22374 3752 22380
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3068 22066 3280 22094
rect 3068 21350 3096 22066
rect 3620 21554 3648 22170
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 2872 20800 2924 20806
rect 2872 20742 2924 20748
rect 3068 20398 3096 21286
rect 3620 20942 3648 21490
rect 3516 20936 3568 20942
rect 3516 20878 3568 20884
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 3528 20754 3556 20878
rect 3528 20726 3648 20754
rect 3620 20466 3648 20726
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 2872 20392 2924 20398
rect 2872 20334 2924 20340
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2424 20058 2452 20198
rect 2884 20058 2912 20334
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 3068 19922 3096 20334
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2976 19446 3004 19654
rect 2964 19440 3016 19446
rect 2964 19382 3016 19388
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2136 17876 2188 17882
rect 2136 17818 2188 17824
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 16574 1992 17478
rect 1872 16546 1992 16574
rect 2136 16584 2188 16590
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1400 16244 1452 16250
rect 1400 16186 1452 16192
rect 1412 16046 1440 16186
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 938 15736 994 15745
rect 938 15671 940 15680
rect 992 15671 994 15680
rect 940 15642 992 15648
rect 1412 14414 1440 15982
rect 1780 15502 1808 16390
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 13394 1440 14350
rect 1676 14340 1728 14346
rect 1676 14282 1728 14288
rect 1688 14074 1716 14282
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1504 13705 1532 13806
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 1400 13388 1452 13394
rect 1400 13330 1452 13336
rect 1412 12850 1440 13330
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 12442 1716 12718
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11665 980 11698
rect 938 11656 994 11665
rect 938 11591 994 11600
rect 1676 11076 1728 11082
rect 1676 11018 1728 11024
rect 1688 10810 1716 11018
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 938 8936 994 8945
rect 938 8871 940 8880
rect 992 8871 994 8880
rect 940 8842 992 8848
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 6905 1532 7346
rect 1872 6914 1900 16546
rect 2516 16574 2544 18022
rect 2136 16526 2188 16532
rect 2424 16546 2544 16574
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 16182 1992 16390
rect 1952 16176 2004 16182
rect 1952 16118 2004 16124
rect 2148 16046 2176 16526
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 1490 6896 1546 6905
rect 1872 6886 1992 6914
rect 1490 6831 1546 6840
rect 940 4548 992 4554
rect 940 4490 992 4496
rect 952 4185 980 4490
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 1964 3058 1992 6886
rect 2424 3058 2452 16546
rect 2976 16250 3004 18022
rect 3068 17066 3096 19858
rect 3160 19242 3188 20402
rect 3620 19378 3648 20402
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 3160 18698 3188 19178
rect 3148 18692 3200 18698
rect 3148 18634 3200 18640
rect 3516 18080 3568 18086
rect 3516 18022 3568 18028
rect 3528 17746 3556 18022
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3436 17338 3464 17614
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3056 17060 3108 17066
rect 3056 17002 3108 17008
rect 3068 16658 3096 17002
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 3068 14940 3096 16594
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3160 15910 3188 16390
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3252 15026 3280 17138
rect 3620 16794 3648 19314
rect 3712 18154 3740 22374
rect 3896 21962 3924 22578
rect 4080 22030 4108 22578
rect 4172 22438 4200 23258
rect 4436 23112 4488 23118
rect 4436 23054 4488 23060
rect 4448 22778 4476 23054
rect 4528 23044 4580 23050
rect 4528 22986 4580 22992
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 4540 22710 4568 22986
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4528 22704 4580 22710
rect 4528 22646 4580 22652
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 3884 21956 3936 21962
rect 3884 21898 3936 21904
rect 3896 20602 3924 21898
rect 4080 21010 4108 21966
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 4356 21690 4384 21830
rect 4344 21684 4396 21690
rect 4632 21672 4660 22918
rect 4724 22642 4752 24160
rect 4816 23322 4844 24686
rect 5632 24608 5684 24614
rect 5632 24550 5684 24556
rect 5644 24274 5672 24550
rect 5632 24268 5684 24274
rect 5632 24210 5684 24216
rect 5632 23724 5684 23730
rect 5632 23666 5684 23672
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 4896 23112 4948 23118
rect 4894 23080 4896 23089
rect 4948 23080 4950 23089
rect 5276 23050 5304 23462
rect 5644 23322 5672 23666
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 5356 23248 5408 23254
rect 5356 23190 5408 23196
rect 5368 23050 5396 23190
rect 4894 23015 4950 23024
rect 5264 23044 5316 23050
rect 5264 22986 5316 22992
rect 5356 23044 5408 23050
rect 5356 22986 5408 22992
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 4712 22636 4764 22642
rect 4712 22578 4764 22584
rect 4712 21684 4764 21690
rect 4632 21644 4712 21672
rect 4344 21626 4396 21632
rect 4712 21626 4764 21632
rect 4620 21412 4672 21418
rect 4620 21354 4672 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21146 4660 21354
rect 4620 21140 4672 21146
rect 4620 21082 4672 21088
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3884 20596 3936 20602
rect 3884 20538 3936 20544
rect 3988 20466 4016 20878
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3792 20324 3844 20330
rect 3792 20266 3844 20272
rect 3804 19854 3832 20266
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3896 19446 3924 19790
rect 3988 19718 4016 20198
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3884 19440 3936 19446
rect 3884 19382 3936 19388
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3700 18148 3752 18154
rect 3700 18090 3752 18096
rect 3712 17678 3740 18090
rect 3988 17746 4016 19246
rect 4080 18834 4108 20742
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4620 19780 4672 19786
rect 4724 19768 4752 21626
rect 4816 19922 4844 22646
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 4908 21434 4936 22510
rect 5184 21622 5212 22578
rect 5368 22574 5396 22986
rect 5644 22778 5672 23258
rect 5828 23254 5856 24890
rect 6012 24886 6040 26182
rect 6932 26042 6960 26182
rect 6920 26036 6972 26042
rect 6920 25978 6972 25984
rect 6000 24880 6052 24886
rect 6000 24822 6052 24828
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 5920 23866 5948 24754
rect 6012 24138 6040 24822
rect 7116 24614 7144 29056
rect 7196 28484 7248 28490
rect 7196 28426 7248 28432
rect 7208 28150 7236 28426
rect 7196 28144 7248 28150
rect 7196 28086 7248 28092
rect 7208 27062 7236 28086
rect 7484 28014 7512 30738
rect 7840 30592 7892 30598
rect 7668 30540 7840 30546
rect 7668 30534 7892 30540
rect 7668 30518 7880 30534
rect 7668 30394 7696 30518
rect 7656 30388 7708 30394
rect 7656 30330 7708 30336
rect 7748 30388 7800 30394
rect 7748 30330 7800 30336
rect 7760 30258 7788 30330
rect 7944 30258 7972 31776
rect 8116 31758 8168 31764
rect 8024 30592 8076 30598
rect 8024 30534 8076 30540
rect 8036 30394 8064 30534
rect 8024 30388 8076 30394
rect 8024 30330 8076 30336
rect 7748 30252 7800 30258
rect 7748 30194 7800 30200
rect 7932 30252 7984 30258
rect 7932 30194 7984 30200
rect 7944 30054 7972 30194
rect 7932 30048 7984 30054
rect 7932 29990 7984 29996
rect 7944 29170 7972 29990
rect 7932 29164 7984 29170
rect 7932 29106 7984 29112
rect 8128 28490 8156 31758
rect 8220 28506 8248 32846
rect 8312 32366 8340 33458
rect 8588 32910 8616 38286
rect 9048 36174 9076 38286
rect 9588 38276 9640 38282
rect 9588 38218 9640 38224
rect 10232 38276 10284 38282
rect 10232 38218 10284 38224
rect 11060 38276 11112 38282
rect 11060 38218 11112 38224
rect 9600 38010 9628 38218
rect 9588 38004 9640 38010
rect 9588 37946 9640 37952
rect 9508 37466 9628 37482
rect 9508 37460 9640 37466
rect 9508 37454 9588 37460
rect 9508 36718 9536 37454
rect 9588 37402 9640 37408
rect 9588 37324 9640 37330
rect 9588 37266 9640 37272
rect 9600 36854 9628 37266
rect 10244 37262 10272 38218
rect 10692 37936 10744 37942
rect 10692 37878 10744 37884
rect 10232 37256 10284 37262
rect 10232 37198 10284 37204
rect 9588 36848 9640 36854
rect 9588 36790 9640 36796
rect 9496 36712 9548 36718
rect 9496 36654 9548 36660
rect 9864 36712 9916 36718
rect 9864 36654 9916 36660
rect 9036 36168 9088 36174
rect 9036 36110 9088 36116
rect 9048 35894 9076 36110
rect 9404 36032 9456 36038
rect 9404 35974 9456 35980
rect 9416 35894 9444 35974
rect 9048 35866 9168 35894
rect 8668 34944 8720 34950
rect 8668 34886 8720 34892
rect 8680 34474 8708 34886
rect 8852 34536 8904 34542
rect 8852 34478 8904 34484
rect 8668 34468 8720 34474
rect 8668 34410 8720 34416
rect 8864 34406 8892 34478
rect 8852 34400 8904 34406
rect 8852 34342 8904 34348
rect 8668 33856 8720 33862
rect 8668 33798 8720 33804
rect 8680 33658 8708 33798
rect 8668 33652 8720 33658
rect 8668 33594 8720 33600
rect 8864 32994 8892 34342
rect 9048 34066 9076 35866
rect 9140 35834 9168 35866
rect 9232 35866 9444 35894
rect 9128 35828 9180 35834
rect 9128 35770 9180 35776
rect 9232 35698 9260 35866
rect 9220 35692 9272 35698
rect 9220 35634 9272 35640
rect 9508 35630 9536 36654
rect 9772 36168 9824 36174
rect 9772 36110 9824 36116
rect 9588 36032 9640 36038
rect 9588 35974 9640 35980
rect 9600 35766 9628 35974
rect 9588 35760 9640 35766
rect 9588 35702 9640 35708
rect 9496 35624 9548 35630
rect 9496 35566 9548 35572
rect 9784 35290 9812 36110
rect 9876 35894 9904 36654
rect 10244 36174 10272 37198
rect 10600 37120 10652 37126
rect 10600 37062 10652 37068
rect 10612 36854 10640 37062
rect 10704 36922 10732 37878
rect 10784 37800 10836 37806
rect 10784 37742 10836 37748
rect 10692 36916 10744 36922
rect 10692 36858 10744 36864
rect 10600 36848 10652 36854
rect 10600 36790 10652 36796
rect 10612 36174 10640 36790
rect 10232 36168 10284 36174
rect 10232 36110 10284 36116
rect 10600 36168 10652 36174
rect 10600 36110 10652 36116
rect 9876 35866 9996 35894
rect 9772 35284 9824 35290
rect 9772 35226 9824 35232
rect 9864 35216 9916 35222
rect 9784 35164 9864 35170
rect 9784 35158 9916 35164
rect 9784 35142 9904 35158
rect 9036 34060 9088 34066
rect 9036 34002 9088 34008
rect 8944 33856 8996 33862
rect 8944 33798 8996 33804
rect 8956 33114 8984 33798
rect 8944 33108 8996 33114
rect 8944 33050 8996 33056
rect 8864 32966 8984 32994
rect 8576 32904 8628 32910
rect 8576 32846 8628 32852
rect 8852 32768 8904 32774
rect 8852 32710 8904 32716
rect 8300 32360 8352 32366
rect 8300 32302 8352 32308
rect 8576 32020 8628 32026
rect 8576 31962 8628 31968
rect 8484 31816 8536 31822
rect 8484 31758 8536 31764
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 8312 31482 8340 31622
rect 8300 31476 8352 31482
rect 8300 31418 8352 31424
rect 8392 31408 8444 31414
rect 8392 31350 8444 31356
rect 8404 30938 8432 31350
rect 8496 30938 8524 31758
rect 8392 30932 8444 30938
rect 8392 30874 8444 30880
rect 8484 30932 8536 30938
rect 8484 30874 8536 30880
rect 8588 30258 8616 31962
rect 8864 31822 8892 32710
rect 8852 31816 8904 31822
rect 8852 31758 8904 31764
rect 8576 30252 8628 30258
rect 8576 30194 8628 30200
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 8312 29306 8340 29582
rect 8392 29572 8444 29578
rect 8392 29514 8444 29520
rect 8300 29300 8352 29306
rect 8300 29242 8352 29248
rect 8298 29200 8354 29209
rect 8404 29186 8432 29514
rect 8354 29158 8432 29186
rect 8298 29135 8354 29144
rect 8588 28994 8616 30194
rect 8588 28966 8800 28994
rect 8392 28960 8444 28966
rect 8484 28960 8536 28966
rect 8444 28920 8484 28948
rect 8392 28902 8444 28908
rect 8484 28902 8536 28908
rect 8496 28762 8524 28902
rect 8484 28756 8536 28762
rect 8484 28698 8536 28704
rect 8116 28484 8168 28490
rect 8220 28478 8340 28506
rect 8116 28426 8168 28432
rect 7932 28416 7984 28422
rect 7932 28358 7984 28364
rect 7944 28150 7972 28358
rect 7932 28144 7984 28150
rect 8312 28098 8340 28478
rect 7932 28086 7984 28092
rect 8220 28070 8340 28098
rect 7472 28008 7524 28014
rect 7472 27950 7524 27956
rect 7196 27056 7248 27062
rect 7196 26998 7248 27004
rect 7380 27056 7432 27062
rect 7380 26998 7432 27004
rect 7392 26790 7420 26998
rect 7484 26926 7512 27950
rect 7564 27328 7616 27334
rect 7564 27270 7616 27276
rect 7472 26920 7524 26926
rect 7472 26862 7524 26868
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7288 26444 7340 26450
rect 7576 26432 7604 27270
rect 7340 26404 7604 26432
rect 7288 26386 7340 26392
rect 7576 25294 7604 26404
rect 7840 26444 7892 26450
rect 8116 26444 8168 26450
rect 7892 26404 8116 26432
rect 7840 26386 7892 26392
rect 8116 26386 8168 26392
rect 7840 26240 7892 26246
rect 8116 26240 8168 26246
rect 7892 26200 8116 26228
rect 7840 26182 7892 26188
rect 8116 26182 8168 26188
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 7300 24750 7328 25094
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7944 24410 7972 24686
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 6000 24132 6052 24138
rect 6000 24074 6052 24080
rect 5908 23860 5960 23866
rect 5908 23802 5960 23808
rect 6012 23594 6040 24074
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6932 23866 6960 24006
rect 6920 23860 6972 23866
rect 6920 23802 6972 23808
rect 7288 23860 7340 23866
rect 7288 23802 7340 23808
rect 6000 23588 6052 23594
rect 6000 23530 6052 23536
rect 6550 23352 6606 23361
rect 6550 23287 6606 23296
rect 5816 23248 5868 23254
rect 5816 23190 5868 23196
rect 5828 23100 5856 23190
rect 6564 23186 6592 23287
rect 6552 23180 6604 23186
rect 6552 23122 6604 23128
rect 5908 23112 5960 23118
rect 5828 23072 5908 23100
rect 6932 23100 6960 23802
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 7024 23322 7052 23666
rect 7300 23594 7328 23802
rect 7288 23588 7340 23594
rect 7288 23530 7340 23536
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7012 23112 7064 23118
rect 6932 23072 7012 23100
rect 5908 23054 5960 23060
rect 7012 23054 7064 23060
rect 5632 22772 5684 22778
rect 5632 22714 5684 22720
rect 5920 22710 5948 23054
rect 6000 22976 6052 22982
rect 6000 22918 6052 22924
rect 5908 22704 5960 22710
rect 5908 22646 5960 22652
rect 5356 22568 5408 22574
rect 5356 22510 5408 22516
rect 6012 22166 6040 22918
rect 7024 22778 7052 23054
rect 7208 23050 7236 23258
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 7012 22772 7064 22778
rect 7012 22714 7064 22720
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6276 22500 6328 22506
rect 6276 22442 6328 22448
rect 6184 22432 6236 22438
rect 6184 22374 6236 22380
rect 6000 22160 6052 22166
rect 6000 22102 6052 22108
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 5172 21616 5224 21622
rect 5172 21558 5224 21564
rect 5828 21554 5856 21830
rect 6196 21554 6224 22374
rect 6288 22166 6316 22442
rect 6276 22160 6328 22166
rect 6276 22102 6328 22108
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 4908 21418 5120 21434
rect 4908 21412 5132 21418
rect 4908 21406 5080 21412
rect 5080 21354 5132 21360
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 4672 19740 4752 19768
rect 4620 19722 4672 19728
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4080 18222 4108 18770
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4264 18426 4292 18566
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3700 17672 3752 17678
rect 3700 17614 3752 17620
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3620 16250 3648 16730
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3148 14952 3200 14958
rect 3068 14912 3148 14940
rect 3148 14894 3200 14900
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2516 14074 2544 14758
rect 2964 14340 3016 14346
rect 2964 14282 3016 14288
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2976 13190 3004 14282
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2976 12850 3004 13126
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2976 11082 3004 12786
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3068 12306 3096 12582
rect 3160 12434 3188 14894
rect 3252 14618 3280 14962
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14618 3648 14758
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3712 14482 3740 17614
rect 4080 17270 4108 18158
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 4264 17338 4292 17546
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3160 12406 3280 12434
rect 3252 12306 3280 12406
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 3148 12164 3200 12170
rect 3148 12106 3200 12112
rect 3160 11354 3188 12106
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 3160 10674 3188 11290
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10062 3188 10610
rect 3252 10470 3280 12242
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3344 10062 3372 13262
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11354 3464 12038
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3436 10606 3464 11290
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3160 9722 3188 9862
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3238 9616 3294 9625
rect 3238 9551 3240 9560
rect 3292 9551 3294 9560
rect 3240 9522 3292 9528
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 9178 3004 9318
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3344 8974 3372 9998
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 7478 3004 8230
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 3620 7342 3648 11494
rect 3712 9586 3740 14418
rect 3804 13326 3832 17070
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16776 4660 19722
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4816 18970 4844 19246
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4264 16748 4660 16776
rect 3976 16584 4028 16590
rect 4160 16584 4212 16590
rect 3976 16526 4028 16532
rect 4080 16544 4160 16572
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15502 3924 15846
rect 3988 15706 4016 16526
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 4080 15586 4108 16544
rect 4160 16526 4212 16532
rect 4264 16522 4292 16748
rect 4436 16652 4488 16658
rect 4488 16612 4568 16640
rect 4436 16594 4488 16600
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 4540 16402 4568 16612
rect 4540 16374 4752 16402
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15638 4660 16186
rect 4724 15706 4752 16374
rect 4816 16182 4844 17206
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4620 15632 4672 15638
rect 4080 15558 4292 15586
rect 4620 15574 4672 15580
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 3988 15026 4016 15438
rect 4172 15094 4200 15438
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 4264 14958 4292 15558
rect 4632 15094 4660 15574
rect 4816 15502 4844 16118
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3896 12782 3924 14758
rect 4080 14618 4108 14826
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4632 14414 4660 15030
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 3988 13002 4016 13194
rect 3988 12986 4108 13002
rect 4632 12986 4660 13194
rect 3976 12980 4108 12986
rect 4028 12974 4108 12980
rect 3976 12922 4028 12928
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3804 12442 3832 12650
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3896 11286 3924 12718
rect 3988 12322 4016 12786
rect 4080 12442 4108 12974
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4724 12850 4752 14962
rect 4436 12844 4488 12850
rect 4712 12844 4764 12850
rect 4488 12804 4660 12832
rect 4436 12786 4488 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12442 4660 12804
rect 4712 12786 4764 12792
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 3988 12306 4108 12322
rect 3988 12300 4120 12306
rect 3988 12294 4068 12300
rect 4068 12242 4120 12248
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10810 3832 10950
rect 3896 10810 3924 11018
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3896 8922 3924 10746
rect 4080 10606 4108 11154
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10742 4292 10950
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3988 9110 4016 9318
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3896 8894 4016 8922
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3896 4622 3924 8774
rect 3988 7410 4016 8894
rect 4080 8362 4108 10542
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4724 10266 4752 10542
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4158 9072 4214 9081
rect 4724 9042 4752 9318
rect 4158 9007 4214 9016
rect 4712 9036 4764 9042
rect 4172 8974 4200 9007
rect 4712 8978 4764 8984
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4724 8498 4752 8842
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7546 4660 8230
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6866 4660 7482
rect 4724 7342 4752 8434
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 4540 6458 4568 6666
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 2228 2848 2280 2854
rect 2228 2790 2280 2796
rect 1780 2446 1808 2790
rect 2240 2446 2268 2790
rect 4908 2774 4936 21286
rect 5092 19718 5120 21354
rect 5736 21185 5764 21490
rect 5722 21176 5778 21185
rect 5722 21111 5778 21120
rect 5630 20904 5686 20913
rect 5630 20839 5632 20848
rect 5684 20839 5686 20848
rect 5632 20810 5684 20816
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5092 19514 5120 19654
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 5184 18766 5212 19654
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5460 17746 5488 19314
rect 5828 18698 5856 21490
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5920 19514 5948 19790
rect 5908 19508 5960 19514
rect 5908 19450 5960 19456
rect 5920 18834 5948 19450
rect 5998 18864 6054 18873
rect 5908 18828 5960 18834
rect 5998 18799 6054 18808
rect 5908 18770 5960 18776
rect 6012 18766 6040 18799
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 5632 18692 5684 18698
rect 5632 18634 5684 18640
rect 5816 18692 5868 18698
rect 5816 18634 5868 18640
rect 5644 17882 5672 18634
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5632 17876 5684 17882
rect 5632 17818 5684 17824
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 5000 16250 5028 17070
rect 5460 16250 5488 17682
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5736 17338 5764 17478
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5920 16522 5948 18158
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6196 17542 6224 18022
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6104 16794 6132 16934
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 5908 16516 5960 16522
rect 5908 16458 5960 16464
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5920 16046 5948 16458
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5908 16040 5960 16046
rect 5908 15982 5960 15988
rect 5644 15706 5672 15982
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 6196 15570 6224 17478
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5460 15162 5488 15302
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5552 9654 5580 13806
rect 5644 13394 5672 14350
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5920 14074 5948 14282
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6288 13394 6316 22102
rect 6932 21894 6960 22578
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 6932 21622 6960 21830
rect 7300 21622 7328 23530
rect 7746 23352 7802 23361
rect 7746 23287 7802 23296
rect 7380 23044 7432 23050
rect 7380 22986 7432 22992
rect 7564 23044 7616 23050
rect 7564 22986 7616 22992
rect 7392 22710 7420 22986
rect 7380 22704 7432 22710
rect 7380 22646 7432 22652
rect 6920 21616 6972 21622
rect 6920 21558 6972 21564
rect 7288 21616 7340 21622
rect 7288 21558 7340 21564
rect 6828 21480 6880 21486
rect 6828 21422 6880 21428
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6656 19854 6684 21286
rect 6840 21146 6868 21422
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 6932 20942 6960 21558
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6564 19514 6592 19790
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 6564 18630 6592 19450
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 6656 18222 6684 19790
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 6932 19514 6960 19722
rect 7208 19514 7236 20198
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 7196 19508 7248 19514
rect 7196 19450 7248 19456
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6748 18290 6776 18566
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6932 17610 6960 17818
rect 6368 17604 6420 17610
rect 6368 17546 6420 17552
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6380 17338 6408 17546
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6932 15434 6960 17546
rect 7392 17542 7420 20334
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7208 17134 7236 17478
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5828 12442 5856 12786
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 6288 12306 6316 13330
rect 6380 12850 6408 15370
rect 6472 15162 6500 15370
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6932 14346 6960 15370
rect 7208 14958 7236 17070
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6932 13394 6960 14282
rect 7208 13870 7236 14894
rect 7484 14618 7512 19994
rect 7576 19718 7604 22986
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 7668 22710 7696 22918
rect 7656 22704 7708 22710
rect 7656 22646 7708 22652
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7760 17882 7788 23287
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7760 17338 7788 17818
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7576 15706 7604 17002
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7576 15162 7604 15642
rect 7852 15502 7880 24346
rect 8022 23080 8078 23089
rect 7932 23044 7984 23050
rect 8022 23015 8078 23024
rect 7932 22986 7984 22992
rect 7944 22710 7972 22986
rect 7932 22704 7984 22710
rect 7932 22646 7984 22652
rect 7932 21004 7984 21010
rect 7932 20946 7984 20952
rect 7944 20398 7972 20946
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7932 19984 7984 19990
rect 7932 19926 7984 19932
rect 7944 19417 7972 19926
rect 7930 19408 7986 19417
rect 7930 19343 7986 19352
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 7944 17882 7972 18158
rect 7932 17876 7984 17882
rect 7932 17818 7984 17824
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7484 14006 7512 14554
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7208 13394 7236 13806
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6564 12986 6592 13126
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6932 12918 6960 13330
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 7208 12434 7236 13330
rect 8036 13190 8064 23015
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 8128 21894 8156 22578
rect 8116 21888 8168 21894
rect 8116 21830 8168 21836
rect 8128 21350 8156 21830
rect 8116 21344 8168 21350
rect 8116 21286 8168 21292
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 8128 14890 8156 19994
rect 8220 19514 8248 28070
rect 8300 28008 8352 28014
rect 8300 27950 8352 27956
rect 8312 27674 8340 27950
rect 8300 27668 8352 27674
rect 8300 27610 8352 27616
rect 8392 26920 8444 26926
rect 8392 26862 8444 26868
rect 8404 26382 8432 26862
rect 8772 26450 8800 28966
rect 8760 26444 8812 26450
rect 8760 26386 8812 26392
rect 8392 26376 8444 26382
rect 8392 26318 8444 26324
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 8496 21894 8524 26250
rect 8668 26240 8720 26246
rect 8668 26182 8720 26188
rect 8680 25838 8708 26182
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8772 22642 8800 26386
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8864 21690 8892 31758
rect 8956 31482 8984 32966
rect 9048 31890 9076 34002
rect 9588 33924 9640 33930
rect 9588 33866 9640 33872
rect 9404 33856 9456 33862
rect 9404 33798 9456 33804
rect 9416 33658 9444 33798
rect 9404 33652 9456 33658
rect 9404 33594 9456 33600
rect 9600 33454 9628 33866
rect 9588 33448 9640 33454
rect 9588 33390 9640 33396
rect 9784 33114 9812 35142
rect 9864 34400 9916 34406
rect 9968 34388 9996 35866
rect 10244 35850 10272 36110
rect 10244 35822 10364 35850
rect 10244 35766 10272 35822
rect 10232 35760 10284 35766
rect 10232 35702 10284 35708
rect 9916 34360 9996 34388
rect 9864 34342 9916 34348
rect 9864 33992 9916 33998
rect 9864 33934 9916 33940
rect 9876 33114 9904 33934
rect 10336 33522 10364 35822
rect 10324 33516 10376 33522
rect 10324 33458 10376 33464
rect 9772 33108 9824 33114
rect 9772 33050 9824 33056
rect 9864 33108 9916 33114
rect 9864 33050 9916 33056
rect 9784 32774 9812 33050
rect 9772 32768 9824 32774
rect 9772 32710 9824 32716
rect 9036 31884 9088 31890
rect 9036 31826 9088 31832
rect 8944 31476 8996 31482
rect 8944 31418 8996 31424
rect 9048 29510 9076 31826
rect 10336 31754 10364 33458
rect 10600 33312 10652 33318
rect 10600 33254 10652 33260
rect 10612 32910 10640 33254
rect 10600 32904 10652 32910
rect 10600 32846 10652 32852
rect 10508 32768 10560 32774
rect 10508 32710 10560 32716
rect 9772 31748 9824 31754
rect 9772 31690 9824 31696
rect 10324 31748 10376 31754
rect 10324 31690 10376 31696
rect 9784 31482 9812 31690
rect 10520 31482 10548 32710
rect 10704 31754 10732 36858
rect 10796 35222 10824 37742
rect 11072 37466 11100 38218
rect 11348 37874 11376 38286
rect 11888 38208 11940 38214
rect 11888 38150 11940 38156
rect 11900 37942 11928 38150
rect 12084 38010 12112 38898
rect 12360 38010 12388 38966
rect 20088 38962 20116 40854
rect 21914 40762 21970 41562
rect 24490 40762 24546 41562
rect 26422 40762 26478 41562
rect 28354 40762 28410 41562
rect 30930 40762 30986 41562
rect 32862 40882 32918 41562
rect 32862 40854 33088 40882
rect 32862 40762 32918 40854
rect 21928 39098 21956 40762
rect 26436 39098 26464 40762
rect 21916 39092 21968 39098
rect 21916 39034 21968 39040
rect 26424 39092 26476 39098
rect 26424 39034 26476 39040
rect 30944 39030 30972 40762
rect 33060 39794 33088 40854
rect 35438 40762 35494 41562
rect 37370 40762 37426 41562
rect 39302 40762 39358 41562
rect 33060 39766 33180 39794
rect 33152 39098 33180 39766
rect 35452 39098 35480 40762
rect 33140 39092 33192 39098
rect 33140 39034 33192 39040
rect 35440 39092 35492 39098
rect 35440 39034 35492 39040
rect 30932 39024 30984 39030
rect 20350 38992 20406 39001
rect 12440 38956 12492 38962
rect 12440 38898 12492 38904
rect 17960 38956 18012 38962
rect 17960 38898 18012 38904
rect 19432 38956 19484 38962
rect 19432 38898 19484 38904
rect 20076 38956 20128 38962
rect 30932 38966 30984 38972
rect 37384 38962 37412 40762
rect 20350 38927 20406 38936
rect 22376 38956 22428 38962
rect 20076 38898 20128 38904
rect 12072 38004 12124 38010
rect 12072 37946 12124 37952
rect 12348 38004 12400 38010
rect 12348 37946 12400 37952
rect 11888 37936 11940 37942
rect 11888 37878 11940 37884
rect 11336 37868 11388 37874
rect 11336 37810 11388 37816
rect 11060 37460 11112 37466
rect 11060 37402 11112 37408
rect 10968 35488 11020 35494
rect 10968 35430 11020 35436
rect 10980 35290 11008 35430
rect 10968 35284 11020 35290
rect 10968 35226 11020 35232
rect 10784 35216 10836 35222
rect 10784 35158 10836 35164
rect 10612 31726 10732 31754
rect 9496 31476 9548 31482
rect 9496 31418 9548 31424
rect 9772 31476 9824 31482
rect 9772 31418 9824 31424
rect 10508 31476 10560 31482
rect 10508 31418 10560 31424
rect 9508 30802 9536 31418
rect 10232 31272 10284 31278
rect 10232 31214 10284 31220
rect 9588 31204 9640 31210
rect 9588 31146 9640 31152
rect 9600 30938 9628 31146
rect 9588 30932 9640 30938
rect 9588 30874 9640 30880
rect 9496 30796 9548 30802
rect 9496 30738 9548 30744
rect 9508 30258 9536 30738
rect 9588 30660 9640 30666
rect 9588 30602 9640 30608
rect 9600 30394 9628 30602
rect 10244 30598 10272 31214
rect 10232 30592 10284 30598
rect 10232 30534 10284 30540
rect 9588 30388 9640 30394
rect 9588 30330 9640 30336
rect 9496 30252 9548 30258
rect 9496 30194 9548 30200
rect 9508 30122 9536 30194
rect 9496 30116 9548 30122
rect 9496 30058 9548 30064
rect 9404 30048 9456 30054
rect 9404 29990 9456 29996
rect 9036 29504 9088 29510
rect 9036 29446 9088 29452
rect 9128 29096 9180 29102
rect 9128 29038 9180 29044
rect 8944 25832 8996 25838
rect 8944 25774 8996 25780
rect 8956 25498 8984 25774
rect 8944 25492 8996 25498
rect 8944 25434 8996 25440
rect 9036 25220 9088 25226
rect 9036 25162 9088 25168
rect 9048 24188 9076 25162
rect 9140 24290 9168 29038
rect 9416 27554 9444 29990
rect 9496 27872 9548 27878
rect 9496 27814 9548 27820
rect 9508 27674 9536 27814
rect 9496 27668 9548 27674
rect 9496 27610 9548 27616
rect 9600 27606 9628 30330
rect 9956 30320 10008 30326
rect 9956 30262 10008 30268
rect 9680 29572 9732 29578
rect 9680 29514 9732 29520
rect 9692 28218 9720 29514
rect 9968 29510 9996 30262
rect 10048 30252 10100 30258
rect 10048 30194 10100 30200
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 9968 28558 9996 29446
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 9680 28212 9732 28218
rect 9680 28154 9732 28160
rect 9772 28076 9824 28082
rect 9772 28018 9824 28024
rect 9680 27872 9732 27878
rect 9680 27814 9732 27820
rect 9692 27674 9720 27814
rect 9680 27668 9732 27674
rect 9680 27610 9732 27616
rect 9588 27600 9640 27606
rect 9416 27526 9536 27554
rect 9588 27542 9640 27548
rect 9220 24948 9272 24954
rect 9220 24890 9272 24896
rect 9232 24410 9260 24890
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9140 24262 9260 24290
rect 9128 24200 9180 24206
rect 9048 24160 9128 24188
rect 9128 24142 9180 24148
rect 9036 24064 9088 24070
rect 9036 24006 9088 24012
rect 9048 23798 9076 24006
rect 9036 23792 9088 23798
rect 9036 23734 9088 23740
rect 9140 23186 9168 24142
rect 9128 23180 9180 23186
rect 9128 23122 9180 23128
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 8300 21412 8352 21418
rect 8300 21354 8352 21360
rect 8312 21146 8340 21354
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8404 19854 8432 20334
rect 8588 20233 8616 21490
rect 8668 20936 8720 20942
rect 8668 20878 8720 20884
rect 8574 20224 8630 20233
rect 8574 20159 8630 20168
rect 8392 19848 8444 19854
rect 8390 19816 8392 19825
rect 8444 19816 8446 19825
rect 8300 19780 8352 19786
rect 8390 19751 8446 19760
rect 8300 19722 8352 19728
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8220 16454 8248 19314
rect 8312 19310 8340 19722
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8312 18358 8340 19246
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8312 17814 8340 18294
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8496 16726 8524 17138
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8312 15162 8340 16594
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12986 8064 13126
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 8128 12434 8156 14826
rect 8312 14006 8340 15098
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8404 13938 8432 14962
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8404 12434 8432 13874
rect 7208 12406 7328 12434
rect 8128 12406 8248 12434
rect 7300 12306 7328 12406
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5644 10742 5672 11154
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5644 8430 5672 10678
rect 5736 10674 5764 11290
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5828 10606 5856 11018
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 10130 5856 10406
rect 5920 10130 5948 11086
rect 6104 10810 6132 11086
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5828 8838 5856 10066
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8480 5856 8774
rect 5920 8634 5948 10066
rect 6104 10062 6132 10746
rect 6748 10674 6776 10950
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 6196 10266 6224 10610
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 10266 6408 10406
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6748 9110 6776 9522
rect 6840 9178 6868 9522
rect 7116 9178 7144 9522
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 7208 8974 7236 10610
rect 7300 9382 7328 12242
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7852 11354 7880 12038
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7484 10674 7512 11086
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7484 10062 7512 10610
rect 7576 10266 7604 11018
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7852 9586 7880 11018
rect 7944 10062 7972 12106
rect 8220 11762 8248 12406
rect 8312 12406 8432 12434
rect 8496 12434 8524 16662
rect 8588 14482 8616 20159
rect 8680 14822 8708 20878
rect 9034 20360 9090 20369
rect 9034 20295 9090 20304
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 8956 19446 8984 19654
rect 9048 19446 9076 20295
rect 8944 19440 8996 19446
rect 8944 19382 8996 19388
rect 9036 19440 9088 19446
rect 9036 19382 9088 19388
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 8772 15162 8800 19314
rect 9140 18086 9168 22714
rect 9232 22094 9260 24262
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9324 23322 9352 23598
rect 9312 23316 9364 23322
rect 9312 23258 9364 23264
rect 9404 23316 9456 23322
rect 9404 23258 9456 23264
rect 9416 23118 9444 23258
rect 9508 23118 9536 27526
rect 9600 26382 9628 27542
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9692 25498 9720 25638
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 9588 25152 9640 25158
rect 9588 25094 9640 25100
rect 9600 24954 9628 25094
rect 9588 24948 9640 24954
rect 9588 24890 9640 24896
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9416 22778 9444 23054
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9692 22234 9720 22986
rect 9680 22228 9732 22234
rect 9680 22170 9732 22176
rect 9232 22066 9352 22094
rect 9324 21690 9352 22066
rect 9784 21894 9812 28018
rect 10060 27996 10088 30194
rect 10140 28008 10192 28014
rect 9968 27968 10140 27996
rect 9864 26852 9916 26858
rect 9864 26794 9916 26800
rect 9876 25362 9904 26794
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 9968 25242 9996 27968
rect 10140 27950 10192 27956
rect 10048 27396 10100 27402
rect 10048 27338 10100 27344
rect 10060 27130 10088 27338
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 10048 25900 10100 25906
rect 10048 25842 10100 25848
rect 9876 25214 9996 25242
rect 9876 24750 9904 25214
rect 9864 24744 9916 24750
rect 9864 24686 9916 24692
rect 9876 24177 9904 24686
rect 9862 24168 9918 24177
rect 9862 24103 9918 24112
rect 9956 23860 10008 23866
rect 10060 23848 10088 25842
rect 10140 25288 10192 25294
rect 10140 25230 10192 25236
rect 10152 24954 10180 25230
rect 10140 24948 10192 24954
rect 10140 24890 10192 24896
rect 10008 23820 10088 23848
rect 9956 23802 10008 23808
rect 10048 23588 10100 23594
rect 10048 23530 10100 23536
rect 10060 23118 10088 23530
rect 10140 23248 10192 23254
rect 10140 23190 10192 23196
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 9876 22778 9904 23054
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 10152 22642 10180 23190
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 10048 22568 10100 22574
rect 10048 22510 10100 22516
rect 10060 22098 10088 22510
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 9678 21584 9734 21593
rect 9678 21519 9680 21528
rect 9732 21519 9734 21528
rect 9680 21490 9732 21496
rect 9784 21146 9812 21830
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9876 21026 9904 21490
rect 9784 20998 9904 21026
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9220 20868 9272 20874
rect 9220 20810 9272 20816
rect 9232 19242 9260 20810
rect 9600 20777 9628 20878
rect 9784 20874 9812 20998
rect 9968 20942 9996 21490
rect 10060 21321 10088 21490
rect 10046 21312 10102 21321
rect 10046 21247 10102 21256
rect 10152 21146 10180 22578
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9864 20868 9916 20874
rect 9864 20810 9916 20816
rect 9586 20768 9642 20777
rect 9586 20703 9642 20712
rect 9784 20534 9812 20810
rect 9772 20528 9824 20534
rect 9772 20470 9824 20476
rect 9494 19952 9550 19961
rect 9494 19887 9550 19896
rect 9508 19854 9536 19887
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9324 19310 9352 19790
rect 9600 19514 9628 19790
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9496 19372 9548 19378
rect 9416 19332 9496 19360
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9220 19236 9272 19242
rect 9220 19178 9272 19184
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 9232 18222 9260 18634
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 8864 16658 8892 18022
rect 9034 17912 9090 17921
rect 8956 17870 9034 17898
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8956 16590 8984 17870
rect 9034 17847 9090 17856
rect 9140 17746 9168 18022
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8956 15178 8984 16526
rect 8760 15156 8812 15162
rect 8956 15150 9076 15178
rect 8760 15098 8812 15104
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8956 14822 8984 14962
rect 9048 14890 9076 15150
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 8668 14816 8720 14822
rect 8944 14816 8996 14822
rect 8720 14776 8892 14804
rect 8668 14758 8720 14764
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8680 14074 8708 14214
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8588 12918 8616 13126
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8496 12406 8616 12434
rect 8312 12238 8340 12406
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8220 11234 8248 11698
rect 8312 11558 8340 12174
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8036 11218 8248 11234
rect 8036 11212 8260 11218
rect 8036 11206 8208 11212
rect 8036 10198 8064 11206
rect 8208 11154 8260 11160
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 8024 10192 8076 10198
rect 8024 10134 8076 10140
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 8128 9586 8156 11018
rect 8312 10470 8340 11494
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8496 10810 8524 11290
rect 8588 11150 8616 12406
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8220 9654 8248 10066
rect 8496 9994 8524 10610
rect 8680 10130 8708 14010
rect 8864 12442 8892 14776
rect 8944 14758 8996 14764
rect 8852 12436 8904 12442
rect 8956 12434 8984 14758
rect 9232 14414 9260 18158
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9048 13530 9076 14350
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 8956 12406 9168 12434
rect 8852 12378 8904 12384
rect 8864 12306 8892 12378
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8772 11898 8800 12174
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8496 9586 8524 9930
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5736 8452 5856 8480
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5552 8090 5580 8366
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5644 7970 5672 8366
rect 5736 8294 5764 8452
rect 5920 8378 5948 8570
rect 6012 8498 6040 8842
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5828 8350 5948 8378
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5828 8090 5856 8350
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5644 7942 5764 7970
rect 5736 7886 5764 7942
rect 5920 7886 5948 8230
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6012 7410 6040 8434
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 7546 6132 7686
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5092 5778 5120 6802
rect 5184 6458 5212 7142
rect 6012 7002 6040 7346
rect 6196 7206 6224 8842
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6380 8294 6408 8434
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7546 6592 7686
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6840 7342 6868 8230
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 6472 5710 6500 6666
rect 6932 5778 6960 7890
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7208 7546 7236 7754
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7484 6254 7512 9386
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 7546 8064 8774
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8220 6798 8248 9386
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8404 8294 8432 8774
rect 8496 8634 8524 8774
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8404 8090 8432 8230
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8220 6322 8248 6734
rect 8496 6662 8524 7754
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5644 5370 5672 5578
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 6932 4146 6960 5714
rect 7392 5370 7420 6054
rect 8220 5914 8248 6054
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8496 5710 8524 6598
rect 8484 5704 8536 5710
rect 8536 5664 8616 5692
rect 8484 5646 8536 5652
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 8220 5234 8248 5510
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8588 4214 8616 5664
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4816 2746 4936 2774
rect 4816 2446 4844 2746
rect 8404 2446 8432 2790
rect 8772 2650 8800 11834
rect 9140 11354 9168 12406
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8864 10674 8892 11222
rect 9140 11150 9168 11290
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 9232 10146 9260 13262
rect 9324 11898 9352 19246
rect 9416 17270 9444 19332
rect 9496 19314 9548 19320
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 9416 16658 9444 17206
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9416 16250 9444 16458
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9508 15162 9536 17274
rect 9600 16998 9628 17478
rect 9692 17270 9720 19790
rect 9784 19718 9812 20470
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9876 17882 9904 20810
rect 9968 19854 9996 20878
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9956 19372 10008 19378
rect 10060 19360 10088 20946
rect 10138 20496 10194 20505
rect 10138 20431 10194 20440
rect 10152 19854 10180 20431
rect 10244 20058 10272 30534
rect 10416 28484 10468 28490
rect 10416 28426 10468 28432
rect 10508 28484 10560 28490
rect 10508 28426 10560 28432
rect 10428 24818 10456 28426
rect 10520 28218 10548 28426
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 10508 25220 10560 25226
rect 10508 25162 10560 25168
rect 10520 24954 10548 25162
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 10612 23254 10640 31726
rect 10968 31476 11020 31482
rect 10968 31418 11020 31424
rect 10980 31278 11008 31418
rect 10968 31272 11020 31278
rect 10968 31214 11020 31220
rect 10692 30116 10744 30122
rect 10692 30058 10744 30064
rect 10704 29850 10732 30058
rect 10692 29844 10744 29850
rect 10692 29786 10744 29792
rect 10704 29306 10732 29786
rect 10692 29300 10744 29306
rect 10692 29242 10744 29248
rect 10980 29102 11008 31214
rect 10968 29096 11020 29102
rect 10968 29038 11020 29044
rect 10980 27878 11008 29038
rect 11072 28490 11100 37402
rect 11348 36174 11376 37810
rect 11704 37800 11756 37806
rect 11702 37768 11704 37777
rect 11756 37768 11758 37777
rect 11702 37703 11758 37712
rect 11520 36576 11572 36582
rect 11520 36518 11572 36524
rect 11532 36174 11560 36518
rect 11704 36304 11756 36310
rect 11704 36246 11756 36252
rect 11336 36168 11388 36174
rect 11336 36110 11388 36116
rect 11520 36168 11572 36174
rect 11520 36110 11572 36116
rect 11152 35760 11204 35766
rect 11152 35702 11204 35708
rect 11060 28484 11112 28490
rect 11060 28426 11112 28432
rect 10968 27872 11020 27878
rect 10968 27814 11020 27820
rect 11072 27470 11100 28426
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 11072 25226 11100 27406
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 10600 23248 10652 23254
rect 10600 23190 10652 23196
rect 11072 23202 11100 25162
rect 11164 23730 11192 35702
rect 11348 35562 11376 36110
rect 11716 35894 11744 36246
rect 11888 36168 11940 36174
rect 11888 36110 11940 36116
rect 12256 36168 12308 36174
rect 12256 36110 12308 36116
rect 11796 36100 11848 36106
rect 11796 36042 11848 36048
rect 11440 35866 11744 35894
rect 11336 35556 11388 35562
rect 11336 35498 11388 35504
rect 11244 26512 11296 26518
rect 11244 26454 11296 26460
rect 11152 23724 11204 23730
rect 11152 23666 11204 23672
rect 11072 23186 11192 23202
rect 11072 23180 11204 23186
rect 11072 23174 11152 23180
rect 11152 23122 11204 23128
rect 11164 23050 11192 23122
rect 11060 23044 11112 23050
rect 11060 22986 11112 22992
rect 11152 23044 11204 23050
rect 11152 22986 11204 22992
rect 11072 22778 11100 22986
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10322 21584 10378 21593
rect 10322 21519 10324 21528
rect 10376 21519 10378 21528
rect 10598 21584 10654 21593
rect 10598 21519 10654 21528
rect 10324 21490 10376 21496
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10008 19332 10088 19360
rect 9956 19314 10008 19320
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9600 15094 9628 16934
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9324 11286 9352 11698
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9416 11234 9444 13670
rect 9508 13190 9536 14894
rect 9586 14376 9642 14385
rect 9586 14311 9588 14320
rect 9640 14311 9642 14320
rect 9588 14282 9640 14288
rect 9586 13696 9642 13705
rect 9586 13631 9642 13640
rect 9600 13394 9628 13631
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9508 12170 9536 13126
rect 9600 12714 9628 13126
rect 9692 12850 9720 16458
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9600 11286 9628 11562
rect 9588 11280 9640 11286
rect 9416 11206 9536 11234
rect 9588 11222 9640 11228
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9416 10810 9444 11086
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9508 10198 9536 11206
rect 8956 10118 9260 10146
rect 9496 10192 9548 10198
rect 9496 10134 9548 10140
rect 8956 10062 8984 10118
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8956 9586 8984 9998
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8864 6118 8892 6326
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8864 5370 8892 6054
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 8956 2514 8984 9522
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9416 7954 9444 8434
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9416 7342 9444 7890
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9508 6798 9536 9862
rect 9692 9466 9720 12786
rect 9784 10130 9812 14758
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9876 12986 9904 14350
rect 9968 13938 9996 19314
rect 10336 18714 10364 21490
rect 10612 20874 10640 21519
rect 10600 20868 10652 20874
rect 10600 20810 10652 20816
rect 10888 18834 10916 21830
rect 11256 21690 11284 26454
rect 11336 22704 11388 22710
rect 11336 22646 11388 22652
rect 11348 22545 11376 22646
rect 11334 22536 11390 22545
rect 11334 22471 11390 22480
rect 11440 22094 11468 35866
rect 11808 35170 11836 36042
rect 11624 35142 11836 35170
rect 11520 34400 11572 34406
rect 11520 34342 11572 34348
rect 11532 33998 11560 34342
rect 11520 33992 11572 33998
rect 11520 33934 11572 33940
rect 11520 32904 11572 32910
rect 11624 32892 11652 35142
rect 11704 34740 11756 34746
rect 11704 34682 11756 34688
rect 11716 34610 11744 34682
rect 11704 34604 11756 34610
rect 11704 34546 11756 34552
rect 11572 32864 11652 32892
rect 11520 32846 11572 32852
rect 11532 30258 11560 32846
rect 11716 32756 11744 34546
rect 11796 34468 11848 34474
rect 11796 34410 11848 34416
rect 11808 33998 11836 34410
rect 11796 33992 11848 33998
rect 11796 33934 11848 33940
rect 11808 33590 11836 33934
rect 11900 33862 11928 36110
rect 11980 36032 12032 36038
rect 11980 35974 12032 35980
rect 11992 34610 12020 35974
rect 12268 34610 12296 36110
rect 11980 34604 12032 34610
rect 11980 34546 12032 34552
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 11888 33856 11940 33862
rect 11888 33798 11940 33804
rect 11796 33584 11848 33590
rect 11796 33526 11848 33532
rect 11796 33312 11848 33318
rect 11796 33254 11848 33260
rect 11808 32910 11836 33254
rect 11796 32904 11848 32910
rect 11796 32846 11848 32852
rect 11796 32768 11848 32774
rect 11716 32728 11796 32756
rect 11796 32710 11848 32716
rect 11612 32224 11664 32230
rect 11612 32166 11664 32172
rect 11624 31958 11652 32166
rect 11612 31952 11664 31958
rect 11612 31894 11664 31900
rect 11612 31680 11664 31686
rect 11612 31622 11664 31628
rect 11624 31346 11652 31622
rect 11612 31340 11664 31346
rect 11612 31282 11664 31288
rect 11624 30870 11652 31282
rect 11612 30864 11664 30870
rect 11612 30806 11664 30812
rect 11704 30728 11756 30734
rect 11704 30670 11756 30676
rect 11716 30258 11744 30670
rect 11808 30410 11836 32710
rect 11900 32434 11928 33798
rect 11992 32842 12020 34546
rect 12072 34060 12124 34066
rect 12072 34002 12124 34008
rect 12084 32881 12112 34002
rect 12070 32872 12126 32881
rect 11980 32836 12032 32842
rect 12070 32807 12072 32816
rect 11980 32778 12032 32784
rect 12124 32807 12126 32816
rect 12072 32778 12124 32784
rect 11888 32428 11940 32434
rect 11888 32370 11940 32376
rect 11900 31346 11928 32370
rect 11992 31414 12020 32778
rect 12268 32298 12296 34546
rect 12348 32768 12400 32774
rect 12348 32710 12400 32716
rect 12360 32570 12388 32710
rect 12348 32564 12400 32570
rect 12348 32506 12400 32512
rect 12256 32292 12308 32298
rect 12256 32234 12308 32240
rect 12268 31754 12296 32234
rect 12176 31726 12296 31754
rect 11980 31408 12032 31414
rect 11980 31350 12032 31356
rect 11888 31340 11940 31346
rect 11888 31282 11940 31288
rect 11808 30382 11928 30410
rect 11900 30258 11928 30382
rect 12176 30258 12204 31726
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 12360 30258 12388 31282
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 11704 30252 11756 30258
rect 11704 30194 11756 30200
rect 11888 30252 11940 30258
rect 11888 30194 11940 30200
rect 12164 30252 12216 30258
rect 12164 30194 12216 30200
rect 12348 30252 12400 30258
rect 12348 30194 12400 30200
rect 11532 28801 11560 30194
rect 11518 28792 11574 28801
rect 11518 28727 11574 28736
rect 11612 27328 11664 27334
rect 11612 27270 11664 27276
rect 11624 27130 11652 27270
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11900 27062 11928 30194
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 11992 28218 12020 28358
rect 11980 28212 12032 28218
rect 11980 28154 12032 28160
rect 11980 28008 12032 28014
rect 11980 27950 12032 27956
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 11992 27538 12020 27950
rect 12084 27878 12112 27950
rect 12072 27872 12124 27878
rect 12072 27814 12124 27820
rect 11980 27532 12032 27538
rect 11980 27474 12032 27480
rect 11888 27056 11940 27062
rect 11888 26998 11940 27004
rect 11900 26382 11928 26998
rect 11888 26376 11940 26382
rect 11888 26318 11940 26324
rect 12084 25378 12112 27814
rect 12176 27130 12204 30194
rect 12256 30048 12308 30054
rect 12256 29990 12308 29996
rect 12268 29850 12296 29990
rect 12256 29844 12308 29850
rect 12256 29786 12308 29792
rect 12254 28792 12310 28801
rect 12254 28727 12310 28736
rect 12164 27124 12216 27130
rect 12164 27066 12216 27072
rect 12268 26994 12296 28727
rect 12348 27328 12400 27334
rect 12348 27270 12400 27276
rect 12360 26994 12388 27270
rect 12256 26988 12308 26994
rect 12256 26930 12308 26936
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 12268 26586 12296 26930
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 12360 26246 12388 26930
rect 12348 26240 12400 26246
rect 12348 26182 12400 26188
rect 12346 25392 12402 25401
rect 12084 25356 12346 25378
rect 12084 25350 12256 25356
rect 12308 25350 12346 25356
rect 12346 25327 12402 25336
rect 12256 25298 12308 25304
rect 11796 25220 11848 25226
rect 11796 25162 11848 25168
rect 11440 22066 11560 22094
rect 11428 22024 11480 22030
rect 11428 21966 11480 21972
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10152 18686 10364 18714
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10060 17746 10088 18566
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 10152 17338 10180 18686
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10244 15706 10272 18294
rect 10336 17678 10364 18566
rect 10784 18352 10836 18358
rect 10784 18294 10836 18300
rect 10796 18154 10824 18294
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10888 18057 10916 18770
rect 10874 18048 10930 18057
rect 10874 17983 10930 17992
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10336 17270 10364 17614
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10244 14482 10272 14758
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 10152 13326 10180 13942
rect 10336 13530 10364 15982
rect 10428 13530 10456 17138
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10140 13320 10192 13326
rect 10060 13280 10140 13308
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9876 11218 9904 12922
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9692 9438 9812 9466
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 7886 9720 9318
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9784 7818 9812 9438
rect 9876 8922 9904 11154
rect 9968 10266 9996 13194
rect 10060 12238 10088 13280
rect 10140 13262 10192 13268
rect 10230 13016 10286 13025
rect 10230 12951 10286 12960
rect 10244 12850 10272 12951
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 9042 10088 9318
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9876 8906 9996 8922
rect 9876 8900 10008 8906
rect 9876 8894 9956 8900
rect 9876 8498 9904 8894
rect 9956 8842 10008 8848
rect 10152 8634 10180 12582
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10244 10606 10272 12174
rect 10336 11694 10364 13466
rect 10428 12986 10456 13466
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10520 12434 10548 17614
rect 10612 17202 10640 17614
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10796 12434 10824 15030
rect 10980 13802 11008 21286
rect 11440 20806 11468 21966
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 11072 17678 11100 19314
rect 11336 19168 11388 19174
rect 11242 19136 11298 19145
rect 11336 19110 11388 19116
rect 11242 19071 11298 19080
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11164 17746 11192 18090
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 11164 17338 11192 17682
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11072 16182 11100 16390
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11256 16046 11284 19071
rect 11348 18630 11376 19110
rect 11440 18834 11468 19654
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11348 18358 11376 18566
rect 11336 18352 11388 18358
rect 11336 18294 11388 18300
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 10428 12406 10548 12434
rect 10704 12406 10824 12434
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10336 11354 10364 11494
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10244 8514 10272 10542
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 10152 8486 10272 8514
rect 9968 7886 9996 8434
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9692 7342 9720 7686
rect 9784 7478 9812 7754
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 5234 9076 6598
rect 9508 6458 9536 6734
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9324 5914 9352 6190
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9416 5710 9444 6326
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5710 9536 6054
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9692 5166 9720 5782
rect 9784 5710 9812 6190
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9140 4282 9168 4966
rect 9692 4282 9720 5102
rect 9784 4622 9812 5646
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9876 5370 9904 5510
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 10060 5234 10088 5510
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9876 4826 9904 5170
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 10152 2650 10180 8486
rect 10428 8430 10456 12406
rect 10704 11762 10732 12406
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10796 11218 10824 11698
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10796 10674 10824 11154
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10612 9042 10640 9590
rect 10704 9586 10732 10134
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10888 9518 10916 11630
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10520 8090 10548 8434
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10888 7750 10916 9454
rect 11072 8378 11100 15642
rect 11334 15600 11390 15609
rect 11244 15564 11296 15570
rect 11334 15535 11390 15544
rect 11244 15506 11296 15512
rect 11256 13530 11284 15506
rect 11348 15502 11376 15535
rect 11336 15496 11388 15502
rect 11388 15456 11468 15484
rect 11532 15473 11560 22066
rect 11808 21894 11836 25162
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 11992 24954 12020 25094
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 12360 24886 12388 25094
rect 12348 24880 12400 24886
rect 12348 24822 12400 24828
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12072 23180 12124 23186
rect 12268 23168 12296 24754
rect 12348 23180 12400 23186
rect 12268 23140 12348 23168
rect 12072 23122 12124 23128
rect 12348 23122 12400 23128
rect 12084 22658 12112 23122
rect 12360 22778 12388 23122
rect 12452 22778 12480 38898
rect 15568 38820 15620 38826
rect 15568 38762 15620 38768
rect 12808 38752 12860 38758
rect 15580 38729 15608 38762
rect 12808 38694 12860 38700
rect 15566 38720 15622 38729
rect 12820 38282 12848 38694
rect 15566 38655 15622 38664
rect 17972 38554 18000 38898
rect 17960 38548 18012 38554
rect 17960 38490 18012 38496
rect 13728 38344 13780 38350
rect 13728 38286 13780 38292
rect 12808 38276 12860 38282
rect 12808 38218 12860 38224
rect 12900 38276 12952 38282
rect 12900 38218 12952 38224
rect 12530 37904 12586 37913
rect 12530 37839 12532 37848
rect 12584 37839 12586 37848
rect 12532 37810 12584 37816
rect 12808 37664 12860 37670
rect 12808 37606 12860 37612
rect 12820 36038 12848 37606
rect 12808 36032 12860 36038
rect 12808 35974 12860 35980
rect 12912 35834 12940 38218
rect 13740 38214 13768 38286
rect 13728 38208 13780 38214
rect 13728 38150 13780 38156
rect 13268 37868 13320 37874
rect 13268 37810 13320 37816
rect 13176 36372 13228 36378
rect 13176 36314 13228 36320
rect 13188 36174 13216 36314
rect 13176 36168 13228 36174
rect 13176 36110 13228 36116
rect 12992 36100 13044 36106
rect 12992 36042 13044 36048
rect 12900 35828 12952 35834
rect 12900 35770 12952 35776
rect 13004 35766 13032 36042
rect 12992 35760 13044 35766
rect 12992 35702 13044 35708
rect 13280 35578 13308 37810
rect 13740 37754 13768 38150
rect 19444 38010 19472 38898
rect 20364 38894 20392 38927
rect 22376 38898 22428 38904
rect 27068 38956 27120 38962
rect 27068 38898 27120 38904
rect 27712 38956 27764 38962
rect 27712 38898 27764 38904
rect 33048 38956 33100 38962
rect 33048 38898 33100 38904
rect 35624 38956 35676 38962
rect 35624 38898 35676 38904
rect 37372 38956 37424 38962
rect 37372 38898 37424 38904
rect 20352 38888 20404 38894
rect 20352 38830 20404 38836
rect 19616 38752 19668 38758
rect 22388 38729 22416 38898
rect 27080 38729 27108 38898
rect 27620 38752 27672 38758
rect 19616 38694 19668 38700
rect 22374 38720 22430 38729
rect 19628 38418 19656 38694
rect 22374 38655 22430 38664
rect 27066 38720 27122 38729
rect 27620 38694 27672 38700
rect 27066 38655 27122 38664
rect 25778 38448 25834 38457
rect 19616 38412 19668 38418
rect 19616 38354 19668 38360
rect 24860 38412 24912 38418
rect 27632 38418 27660 38694
rect 27724 38554 27752 38898
rect 29736 38820 29788 38826
rect 29736 38762 29788 38768
rect 27712 38548 27764 38554
rect 27712 38490 27764 38496
rect 25778 38383 25834 38392
rect 26056 38412 26108 38418
rect 24860 38354 24912 38360
rect 20812 38344 20864 38350
rect 20812 38286 20864 38292
rect 21272 38344 21324 38350
rect 21272 38286 21324 38292
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 15292 38004 15344 38010
rect 15292 37946 15344 37952
rect 16304 38004 16356 38010
rect 16304 37946 16356 37952
rect 19432 38004 19484 38010
rect 19432 37946 19484 37952
rect 14280 37936 14332 37942
rect 14280 37878 14332 37884
rect 13820 37868 13872 37874
rect 13820 37810 13872 37816
rect 13464 37726 13768 37754
rect 13360 35828 13412 35834
rect 13360 35770 13412 35776
rect 13004 35550 13308 35578
rect 12532 35488 12584 35494
rect 12532 35430 12584 35436
rect 12544 34406 12572 35430
rect 12532 34400 12584 34406
rect 12532 34342 12584 34348
rect 12624 33040 12676 33046
rect 12624 32982 12676 32988
rect 12532 31408 12584 31414
rect 12532 31350 12584 31356
rect 12544 28218 12572 31350
rect 12636 29850 12664 32982
rect 13004 31929 13032 35550
rect 13084 34944 13136 34950
rect 13084 34886 13136 34892
rect 12990 31920 13046 31929
rect 12990 31855 13046 31864
rect 12900 31748 12952 31754
rect 12900 31690 12952 31696
rect 12912 31278 12940 31690
rect 12900 31272 12952 31278
rect 12900 31214 12952 31220
rect 12624 29844 12676 29850
rect 12624 29786 12676 29792
rect 12716 29640 12768 29646
rect 12716 29582 12768 29588
rect 12728 29170 12756 29582
rect 12716 29164 12768 29170
rect 12716 29106 12768 29112
rect 12532 28212 12584 28218
rect 12584 28172 12664 28200
rect 12532 28154 12584 28160
rect 12532 27396 12584 27402
rect 12532 27338 12584 27344
rect 12544 26858 12572 27338
rect 12532 26852 12584 26858
rect 12532 26794 12584 26800
rect 12636 26466 12664 28172
rect 12544 26438 12664 26466
rect 12544 25226 12572 26438
rect 12624 26376 12676 26382
rect 12624 26318 12676 26324
rect 12636 25294 12664 26318
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12532 25220 12584 25226
rect 12532 25162 12584 25168
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12544 23662 12572 24550
rect 12728 24274 12756 29106
rect 12898 29064 12954 29073
rect 12898 28999 12900 29008
rect 12952 28999 12954 29008
rect 12900 28970 12952 28976
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12820 25158 12848 26930
rect 12900 26784 12952 26790
rect 12900 26726 12952 26732
rect 12912 26450 12940 26726
rect 12900 26444 12952 26450
rect 12900 26386 12952 26392
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12716 24268 12768 24274
rect 12716 24210 12768 24216
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 12636 23497 12664 24006
rect 12728 23798 12756 24210
rect 12716 23792 12768 23798
rect 12716 23734 12768 23740
rect 13004 23730 13032 31855
rect 13096 29594 13124 34886
rect 13176 34400 13228 34406
rect 13176 34342 13228 34348
rect 13188 34066 13216 34342
rect 13176 34060 13228 34066
rect 13176 34002 13228 34008
rect 13372 33998 13400 35770
rect 13360 33992 13412 33998
rect 13360 33934 13412 33940
rect 13268 33856 13320 33862
rect 13268 33798 13320 33804
rect 13280 33522 13308 33798
rect 13372 33658 13400 33934
rect 13360 33652 13412 33658
rect 13360 33594 13412 33600
rect 13268 33516 13320 33522
rect 13268 33458 13320 33464
rect 13280 31754 13308 33458
rect 13268 31748 13320 31754
rect 13268 31690 13320 31696
rect 13280 30666 13308 31690
rect 13372 31686 13400 33594
rect 13360 31680 13412 31686
rect 13360 31622 13412 31628
rect 13372 30666 13400 31622
rect 13464 31482 13492 37726
rect 13832 36378 13860 37810
rect 14096 37732 14148 37738
rect 14096 37674 14148 37680
rect 13636 36372 13688 36378
rect 13636 36314 13688 36320
rect 13820 36372 13872 36378
rect 13820 36314 13872 36320
rect 13544 35692 13596 35698
rect 13544 35634 13596 35640
rect 13556 33522 13584 35634
rect 13648 35630 13676 36314
rect 14108 36174 14136 37674
rect 14292 36786 14320 37878
rect 14372 37868 14424 37874
rect 14372 37810 14424 37816
rect 14556 37868 14608 37874
rect 14556 37810 14608 37816
rect 14280 36780 14332 36786
rect 14280 36722 14332 36728
rect 14384 36224 14412 37810
rect 14568 36378 14596 37810
rect 14832 36780 14884 36786
rect 14832 36722 14884 36728
rect 14556 36372 14608 36378
rect 14556 36314 14608 36320
rect 14384 36196 14780 36224
rect 14096 36168 14148 36174
rect 14096 36110 14148 36116
rect 14280 36168 14332 36174
rect 14280 36110 14332 36116
rect 14292 35834 14320 36110
rect 14556 36100 14608 36106
rect 14556 36042 14608 36048
rect 14280 35828 14332 35834
rect 14280 35770 14332 35776
rect 13728 35692 13780 35698
rect 13728 35634 13780 35640
rect 13636 35624 13688 35630
rect 13636 35566 13688 35572
rect 13648 34746 13676 35566
rect 13636 34740 13688 34746
rect 13636 34682 13688 34688
rect 13740 33862 13768 35634
rect 14004 34468 14056 34474
rect 14004 34410 14056 34416
rect 13728 33856 13780 33862
rect 13728 33798 13780 33804
rect 13544 33516 13596 33522
rect 13544 33458 13596 33464
rect 13544 32428 13596 32434
rect 13544 32370 13596 32376
rect 13556 32026 13584 32370
rect 13636 32292 13688 32298
rect 13636 32234 13688 32240
rect 13648 32065 13676 32234
rect 13634 32056 13690 32065
rect 13544 32020 13596 32026
rect 13634 31991 13690 32000
rect 13544 31962 13596 31968
rect 13452 31476 13504 31482
rect 13452 31418 13504 31424
rect 13268 30660 13320 30666
rect 13268 30602 13320 30608
rect 13360 30660 13412 30666
rect 13360 30602 13412 30608
rect 13280 29730 13308 30602
rect 13464 30394 13492 31418
rect 13544 31136 13596 31142
rect 13544 31078 13596 31084
rect 13452 30388 13504 30394
rect 13452 30330 13504 30336
rect 13280 29702 13492 29730
rect 13096 29566 13400 29594
rect 13268 29504 13320 29510
rect 13268 29446 13320 29452
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 13188 27470 13216 28018
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 13096 25498 13124 25638
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 13096 25294 13124 25434
rect 13176 25356 13228 25362
rect 13176 25298 13228 25304
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 13188 24886 13216 25298
rect 13176 24880 13228 24886
rect 13176 24822 13228 24828
rect 13176 24608 13228 24614
rect 13176 24550 13228 24556
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12622 23488 12678 23497
rect 12622 23423 12678 23432
rect 12716 23112 12768 23118
rect 12716 23054 12768 23060
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12084 22630 12296 22658
rect 12544 22642 12572 22918
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 11992 22234 12020 22510
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 12176 22098 12204 22510
rect 12164 22092 12216 22098
rect 12164 22034 12216 22040
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 11612 20392 11664 20398
rect 11612 20334 11664 20340
rect 11624 20058 11652 20334
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11624 17746 11652 19994
rect 11716 18442 11744 21830
rect 11808 19990 11836 21830
rect 12176 21486 12204 21830
rect 11980 21480 12032 21486
rect 11980 21422 12032 21428
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 11992 20466 12020 21422
rect 12176 21146 12204 21422
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 12268 20330 12296 22630
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12452 22216 12480 22578
rect 12728 22216 12756 23054
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12452 22188 12756 22216
rect 12452 21554 12480 22188
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12348 21004 12400 21010
rect 12820 20992 12848 22510
rect 12348 20946 12400 20952
rect 12728 20964 12848 20992
rect 12256 20324 12308 20330
rect 12256 20266 12308 20272
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11796 19984 11848 19990
rect 11796 19926 11848 19932
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11808 19514 11836 19654
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11900 19378 11928 20198
rect 12268 19938 12296 20266
rect 11992 19910 12296 19938
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11796 19304 11848 19310
rect 11848 19252 11928 19258
rect 11796 19246 11928 19252
rect 11808 19230 11928 19246
rect 11900 18766 11928 19230
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11716 18414 11836 18442
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11716 17882 11744 18226
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11624 17202 11652 17682
rect 11808 17202 11836 18414
rect 11900 17678 11928 18702
rect 11992 17864 12020 19910
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 12084 19428 12112 19790
rect 12164 19440 12216 19446
rect 12084 19400 12164 19428
rect 12164 19382 12216 19388
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12084 18766 12112 19246
rect 12176 19242 12204 19382
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12164 19236 12216 19242
rect 12164 19178 12216 19184
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12084 18222 12112 18702
rect 12268 18358 12296 19314
rect 12360 18766 12388 20946
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12544 19378 12572 19790
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12360 18290 12388 18702
rect 12544 18698 12572 19314
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12072 18216 12124 18222
rect 12360 18170 12388 18226
rect 12072 18158 12124 18164
rect 12176 18142 12388 18170
rect 11992 17836 12112 17864
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11992 17338 12020 17682
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11808 16998 11836 17138
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11624 15638 11652 15982
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11336 15438 11388 15444
rect 11440 13852 11468 15456
rect 11518 15464 11574 15473
rect 11518 15399 11574 15408
rect 11532 15366 11560 15399
rect 11716 15366 11744 16458
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11440 13824 11652 13852
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11164 12442 11192 13194
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 11256 10606 11284 13466
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11348 11082 11376 11834
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11348 9602 11376 11018
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11440 9722 11468 9998
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11624 9654 11652 13824
rect 11900 13394 11928 15438
rect 11992 14822 12020 16662
rect 12084 16538 12112 17836
rect 12176 17542 12204 18142
rect 12544 17882 12572 18226
rect 12728 18222 12756 20964
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12820 19666 12848 20742
rect 12912 19990 12940 23666
rect 13188 22094 13216 24550
rect 13096 22066 13216 22094
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 12900 19984 12952 19990
rect 12900 19926 12952 19932
rect 12898 19680 12954 19689
rect 12820 19638 12898 19666
rect 12898 19615 12954 19624
rect 12912 19174 12940 19615
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12532 17876 12584 17882
rect 12584 17836 12664 17864
rect 12532 17818 12584 17824
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12360 17542 12388 17614
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12176 17184 12204 17478
rect 12268 17338 12296 17478
rect 12452 17338 12480 17818
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12544 17218 12572 17682
rect 12256 17196 12308 17202
rect 12176 17156 12256 17184
rect 12256 17138 12308 17144
rect 12360 17190 12572 17218
rect 12636 17202 12664 17836
rect 12820 17610 12848 18226
rect 12808 17604 12860 17610
rect 12808 17546 12860 17552
rect 12624 17196 12676 17202
rect 12268 16726 12296 17138
rect 12360 17134 12388 17190
rect 12624 17138 12676 17144
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 12084 16510 12388 16538
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12268 16114 12296 16390
rect 12360 16232 12388 16510
rect 12532 16244 12584 16250
rect 12360 16204 12480 16232
rect 12346 16144 12402 16153
rect 12256 16108 12308 16114
rect 12346 16079 12348 16088
rect 12256 16050 12308 16056
rect 12400 16079 12402 16088
rect 12348 16050 12400 16056
rect 12268 16017 12296 16050
rect 12254 16008 12310 16017
rect 12164 15972 12216 15978
rect 12452 15994 12480 16204
rect 12532 16186 12584 16192
rect 12254 15943 12310 15952
rect 12360 15966 12480 15994
rect 12164 15914 12216 15920
rect 12176 15162 12204 15914
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 12176 14482 12204 15098
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12268 14346 12296 15302
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11900 12850 11928 13330
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11900 11762 11928 12786
rect 11992 12782 12020 14010
rect 12268 13258 12296 14282
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11992 12306 12020 12718
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 12268 11898 12296 13194
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12360 11778 12388 15966
rect 12440 15428 12492 15434
rect 12440 15370 12492 15376
rect 12452 15162 12480 15370
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12544 13734 12572 16186
rect 12820 14958 12848 17546
rect 13004 16182 13032 21830
rect 13096 17882 13124 22066
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 13188 19514 13216 20538
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 12992 16176 13044 16182
rect 12992 16118 13044 16124
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12636 14482 12664 14894
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12544 13326 12572 13670
rect 12636 13394 12664 14418
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12636 12306 12664 13330
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12850 12756 13126
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 11888 11756 11940 11762
rect 11808 11716 11888 11744
rect 11808 10266 11836 11716
rect 11888 11698 11940 11704
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 12084 11750 12388 11778
rect 11992 11354 12020 11698
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11612 9648 11664 9654
rect 11348 9574 11468 9602
rect 11612 9590 11664 9596
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11440 9450 11468 9574
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11348 8634 11376 8910
rect 11440 8906 11468 9386
rect 11624 9178 11652 9590
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11716 8906 11744 9590
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 10980 8350 11100 8378
rect 10980 7886 11008 8350
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 11164 7206 11192 8434
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11532 7342 11560 8026
rect 11808 7478 11836 8434
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11900 7954 11928 8366
rect 12084 7970 12112 11750
rect 12636 11150 12664 12242
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12164 10260 12216 10266
rect 12268 10248 12296 10542
rect 12360 10266 12388 10950
rect 12216 10220 12296 10248
rect 12164 10202 12216 10208
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12176 9450 12204 9862
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12268 8634 12296 10220
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12636 9518 12664 11086
rect 12820 11082 12848 13874
rect 13096 12434 13124 17478
rect 13188 16250 13216 19450
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13004 12406 13124 12434
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12912 11218 12940 11630
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12808 11076 12860 11082
rect 12808 11018 12860 11024
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12162 8528 12218 8537
rect 12162 8463 12218 8472
rect 12176 8362 12204 8463
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12268 8090 12296 8570
rect 12636 8566 12664 9454
rect 13004 8922 13032 12406
rect 13188 12306 13216 12718
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13096 9722 13124 10202
rect 13280 10062 13308 29446
rect 13372 21554 13400 29566
rect 13464 28558 13492 29702
rect 13556 29646 13584 31078
rect 13740 30666 13768 33798
rect 13912 33652 13964 33658
rect 13912 33594 13964 33600
rect 13924 31754 13952 33594
rect 14016 33454 14044 34410
rect 14280 34128 14332 34134
rect 14280 34070 14332 34076
rect 14372 34128 14424 34134
rect 14372 34070 14424 34076
rect 14464 34128 14516 34134
rect 14464 34070 14516 34076
rect 14292 33833 14320 34070
rect 14278 33824 14334 33833
rect 14278 33759 14334 33768
rect 14004 33448 14056 33454
rect 14004 33390 14056 33396
rect 13912 31748 13964 31754
rect 13912 31690 13964 31696
rect 13728 30660 13780 30666
rect 13728 30602 13780 30608
rect 13740 30410 13768 30602
rect 13740 30382 13860 30410
rect 13728 30252 13780 30258
rect 13728 30194 13780 30200
rect 13544 29640 13596 29646
rect 13544 29582 13596 29588
rect 13740 29034 13768 30194
rect 13728 29028 13780 29034
rect 13728 28970 13780 28976
rect 13452 28552 13504 28558
rect 13452 28494 13504 28500
rect 13464 28218 13492 28494
rect 13452 28212 13504 28218
rect 13452 28154 13504 28160
rect 13636 27872 13688 27878
rect 13636 27814 13688 27820
rect 13544 27464 13596 27470
rect 13544 27406 13596 27412
rect 13452 26580 13504 26586
rect 13452 26522 13504 26528
rect 13464 25294 13492 26522
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 13464 23798 13492 25230
rect 13556 24818 13584 27406
rect 13648 26382 13676 27814
rect 13740 27538 13768 28970
rect 13728 27532 13780 27538
rect 13728 27474 13780 27480
rect 13832 27470 13860 30382
rect 13924 29730 13952 31690
rect 14384 30818 14412 34070
rect 14476 33998 14504 34070
rect 14464 33992 14516 33998
rect 14464 33934 14516 33940
rect 14568 33862 14596 36042
rect 14752 33969 14780 36196
rect 14844 36174 14872 36722
rect 15304 36378 15332 37946
rect 16028 37868 16080 37874
rect 16028 37810 16080 37816
rect 16120 37868 16172 37874
rect 16120 37810 16172 37816
rect 16212 37868 16264 37874
rect 16212 37810 16264 37816
rect 16040 37330 16068 37810
rect 15844 37324 15896 37330
rect 15844 37266 15896 37272
rect 16028 37324 16080 37330
rect 16028 37266 16080 37272
rect 15660 36576 15712 36582
rect 15660 36518 15712 36524
rect 15752 36576 15804 36582
rect 15752 36518 15804 36524
rect 15200 36372 15252 36378
rect 15200 36314 15252 36320
rect 15292 36372 15344 36378
rect 15292 36314 15344 36320
rect 14832 36168 14884 36174
rect 14832 36110 14884 36116
rect 14844 34202 14872 36110
rect 15108 36100 15160 36106
rect 15108 36042 15160 36048
rect 15120 35154 15148 36042
rect 15108 35148 15160 35154
rect 15108 35090 15160 35096
rect 14924 34536 14976 34542
rect 14924 34478 14976 34484
rect 14832 34196 14884 34202
rect 14832 34138 14884 34144
rect 14738 33960 14794 33969
rect 14738 33895 14794 33904
rect 14556 33856 14608 33862
rect 14556 33798 14608 33804
rect 14648 33856 14700 33862
rect 14648 33798 14700 33804
rect 14464 31816 14516 31822
rect 14464 31758 14516 31764
rect 14476 30938 14504 31758
rect 14464 30932 14516 30938
rect 14464 30874 14516 30880
rect 14384 30790 14504 30818
rect 14476 30734 14504 30790
rect 14464 30728 14516 30734
rect 14464 30670 14516 30676
rect 14096 30592 14148 30598
rect 14096 30534 14148 30540
rect 14372 30592 14424 30598
rect 14372 30534 14424 30540
rect 13924 29702 14044 29730
rect 13912 29640 13964 29646
rect 13912 29582 13964 29588
rect 13924 28937 13952 29582
rect 13910 28928 13966 28937
rect 13910 28863 13966 28872
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 13636 26376 13688 26382
rect 13924 26364 13952 28863
rect 14016 28218 14044 29702
rect 14108 29646 14136 30534
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 14096 28484 14148 28490
rect 14096 28426 14148 28432
rect 14004 28212 14056 28218
rect 14004 28154 14056 28160
rect 14108 27606 14136 28426
rect 14188 27872 14240 27878
rect 14188 27814 14240 27820
rect 14096 27600 14148 27606
rect 14096 27542 14148 27548
rect 14004 27056 14056 27062
rect 14200 27044 14228 27814
rect 14292 27334 14320 28494
rect 14384 28082 14412 30534
rect 14372 28076 14424 28082
rect 14372 28018 14424 28024
rect 14384 27334 14412 28018
rect 14476 27878 14504 30670
rect 14568 30122 14596 33798
rect 14660 33658 14688 33798
rect 14648 33652 14700 33658
rect 14648 33594 14700 33600
rect 14648 31136 14700 31142
rect 14648 31078 14700 31084
rect 14660 30734 14688 31078
rect 14752 30734 14780 33895
rect 14648 30728 14700 30734
rect 14648 30670 14700 30676
rect 14740 30728 14792 30734
rect 14740 30670 14792 30676
rect 14556 30116 14608 30122
rect 14556 30058 14608 30064
rect 14568 28082 14596 30058
rect 14556 28076 14608 28082
rect 14556 28018 14608 28024
rect 14648 27940 14700 27946
rect 14648 27882 14700 27888
rect 14464 27872 14516 27878
rect 14464 27814 14516 27820
rect 14660 27674 14688 27882
rect 14648 27668 14700 27674
rect 14648 27610 14700 27616
rect 14752 27554 14780 30670
rect 14830 27976 14886 27985
rect 14830 27911 14886 27920
rect 14660 27526 14780 27554
rect 14464 27396 14516 27402
rect 14464 27338 14516 27344
rect 14280 27328 14332 27334
rect 14280 27270 14332 27276
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14056 27016 14228 27044
rect 14004 26998 14056 27004
rect 14292 26976 14320 27270
rect 14372 27056 14424 27062
rect 14372 26998 14424 27004
rect 14108 26948 14320 26976
rect 14004 26376 14056 26382
rect 13924 26336 14004 26364
rect 13636 26318 13688 26324
rect 14004 26318 14056 26324
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13726 24440 13782 24449
rect 13726 24375 13782 24384
rect 13740 24274 13768 24375
rect 13728 24268 13780 24274
rect 13728 24210 13780 24216
rect 13452 23792 13504 23798
rect 13452 23734 13504 23740
rect 13728 23656 13780 23662
rect 13726 23624 13728 23633
rect 13780 23624 13782 23633
rect 13726 23559 13782 23568
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13464 22642 13492 22918
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13740 22030 13768 23559
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13636 21480 13688 21486
rect 13556 21440 13636 21468
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 13464 19718 13492 19926
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13372 19378 13400 19654
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 13372 17746 13400 18634
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13372 15978 13400 17682
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13372 13938 13400 14962
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13372 13394 13400 13874
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13188 9382 13216 9590
rect 13280 9518 13308 9998
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13372 8974 13400 11018
rect 13464 9926 13492 19654
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13360 8968 13412 8974
rect 13004 8894 13216 8922
rect 13360 8910 13412 8916
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 13096 8566 13124 8774
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12360 8248 12480 8276
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12360 7970 12388 8248
rect 11888 7948 11940 7954
rect 12084 7942 12388 7970
rect 11888 7890 11940 7896
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 11796 7472 11848 7478
rect 11796 7414 11848 7420
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 6934 11192 7142
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10244 4622 10272 6258
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10336 5710 10364 5850
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10428 5302 10456 5578
rect 11532 5370 11560 7278
rect 12360 7002 12388 7754
rect 12452 7478 12480 8248
rect 12544 8090 12572 8434
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12452 6338 12480 7414
rect 12820 7002 12848 8230
rect 13004 8090 13032 8434
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13188 7546 13216 8894
rect 13464 8838 13492 9658
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13372 7206 13400 7822
rect 13556 7274 13584 21440
rect 13636 21422 13688 21428
rect 13726 21448 13782 21457
rect 13726 21383 13782 21392
rect 13740 19854 13768 21383
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13648 17542 13676 19722
rect 13726 19544 13782 19553
rect 13726 19479 13782 19488
rect 13740 19446 13768 19479
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13832 18426 13860 25842
rect 14016 24426 14044 26318
rect 14108 24614 14136 26948
rect 14188 26852 14240 26858
rect 14188 26794 14240 26800
rect 14200 25945 14228 26794
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14292 26586 14320 26726
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14384 26466 14412 26998
rect 14292 26450 14412 26466
rect 14280 26444 14412 26450
rect 14332 26438 14412 26444
rect 14280 26386 14332 26392
rect 14186 25936 14242 25945
rect 14186 25871 14242 25880
rect 14188 25220 14240 25226
rect 14188 25162 14240 25168
rect 14200 24954 14228 25162
rect 14188 24948 14240 24954
rect 14188 24890 14240 24896
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14016 24398 14136 24426
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13924 23798 13952 24006
rect 13912 23792 13964 23798
rect 13912 23734 13964 23740
rect 13924 21622 13952 23734
rect 14004 23044 14056 23050
rect 14004 22986 14056 22992
rect 14016 22710 14044 22986
rect 14108 22778 14136 24398
rect 14292 23798 14320 26386
rect 14476 23798 14504 27338
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14568 26466 14596 27270
rect 14660 27062 14688 27526
rect 14648 27056 14700 27062
rect 14648 26998 14700 27004
rect 14738 27024 14794 27033
rect 14738 26959 14740 26968
rect 14792 26959 14794 26968
rect 14740 26930 14792 26936
rect 14648 26920 14700 26926
rect 14648 26862 14700 26868
rect 14660 26586 14688 26862
rect 14648 26580 14700 26586
rect 14648 26522 14700 26528
rect 14568 26438 14688 26466
rect 14556 26308 14608 26314
rect 14556 26250 14608 26256
rect 14568 24886 14596 26250
rect 14660 25838 14688 26438
rect 14648 25832 14700 25838
rect 14648 25774 14700 25780
rect 14556 24880 14608 24886
rect 14556 24822 14608 24828
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14568 24138 14596 24686
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 14280 23792 14332 23798
rect 14278 23760 14280 23769
rect 14464 23792 14516 23798
rect 14332 23760 14334 23769
rect 14188 23724 14240 23730
rect 14464 23734 14516 23740
rect 14278 23695 14334 23704
rect 14188 23666 14240 23672
rect 14200 23322 14228 23666
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 14464 23044 14516 23050
rect 14464 22986 14516 22992
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 14004 22704 14056 22710
rect 14004 22646 14056 22652
rect 14476 22642 14504 22986
rect 14188 22636 14240 22642
rect 14188 22578 14240 22584
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14200 22438 14228 22578
rect 14188 22432 14240 22438
rect 14568 22386 14596 23598
rect 14660 23050 14688 25774
rect 14844 25362 14872 27911
rect 14936 26518 14964 34478
rect 15016 30388 15068 30394
rect 15016 30330 15068 30336
rect 15028 29578 15056 30330
rect 15120 29646 15148 35090
rect 15212 30258 15240 36314
rect 15672 36174 15700 36518
rect 15764 36174 15792 36518
rect 15660 36168 15712 36174
rect 15660 36110 15712 36116
rect 15752 36168 15804 36174
rect 15752 36110 15804 36116
rect 15568 36100 15620 36106
rect 15568 36042 15620 36048
rect 15580 34377 15608 36042
rect 15856 36038 15884 37266
rect 16132 36224 16160 37810
rect 16040 36196 16160 36224
rect 15844 36032 15896 36038
rect 15844 35974 15896 35980
rect 15566 34368 15622 34377
rect 15488 34326 15566 34354
rect 15382 34096 15438 34105
rect 15382 34031 15384 34040
rect 15436 34031 15438 34040
rect 15384 34002 15436 34008
rect 15488 33810 15516 34326
rect 15566 34303 15622 34312
rect 16040 34082 16068 36196
rect 16224 36174 16252 37810
rect 16212 36168 16264 36174
rect 16212 36110 16264 36116
rect 16120 36100 16172 36106
rect 16120 36042 16172 36048
rect 16132 35018 16160 36042
rect 16224 35630 16252 36110
rect 16212 35624 16264 35630
rect 16212 35566 16264 35572
rect 16120 35012 16172 35018
rect 16120 34954 16172 34960
rect 16040 34054 16160 34082
rect 16028 33992 16080 33998
rect 16028 33934 16080 33940
rect 16040 33862 16068 33934
rect 15396 33782 15516 33810
rect 15660 33856 15712 33862
rect 15660 33798 15712 33804
rect 16028 33856 16080 33862
rect 16028 33798 16080 33804
rect 15396 30410 15424 33782
rect 15672 32230 15700 33798
rect 15752 33380 15804 33386
rect 15752 33322 15804 33328
rect 15764 32910 15792 33322
rect 15752 32904 15804 32910
rect 15752 32846 15804 32852
rect 15844 32904 15896 32910
rect 15844 32846 15896 32852
rect 15660 32224 15712 32230
rect 15660 32166 15712 32172
rect 15476 31816 15528 31822
rect 15476 31758 15528 31764
rect 15488 31346 15516 31758
rect 15856 31754 15884 32846
rect 16132 32366 16160 34054
rect 16316 33998 16344 37946
rect 16488 37868 16540 37874
rect 16856 37868 16908 37874
rect 16540 37828 16620 37856
rect 16488 37810 16540 37816
rect 16488 37664 16540 37670
rect 16488 37606 16540 37612
rect 16500 37466 16528 37606
rect 16488 37460 16540 37466
rect 16488 37402 16540 37408
rect 16396 34672 16448 34678
rect 16396 34614 16448 34620
rect 16408 33998 16436 34614
rect 16486 34232 16542 34241
rect 16486 34167 16488 34176
rect 16540 34167 16542 34176
rect 16488 34138 16540 34144
rect 16212 33992 16264 33998
rect 16212 33934 16264 33940
rect 16304 33992 16356 33998
rect 16304 33934 16356 33940
rect 16396 33992 16448 33998
rect 16448 33952 16528 33980
rect 16396 33934 16448 33940
rect 16224 33318 16252 33934
rect 16212 33312 16264 33318
rect 16212 33254 16264 33260
rect 16224 32910 16252 33254
rect 16212 32904 16264 32910
rect 16212 32846 16264 32852
rect 16120 32360 16172 32366
rect 16120 32302 16172 32308
rect 15764 31726 15884 31754
rect 15764 31346 15792 31726
rect 15842 31512 15898 31521
rect 15842 31447 15898 31456
rect 15856 31414 15884 31447
rect 16132 31414 16160 32302
rect 15844 31408 15896 31414
rect 15844 31350 15896 31356
rect 16120 31408 16172 31414
rect 16120 31350 16172 31356
rect 15476 31340 15528 31346
rect 15476 31282 15528 31288
rect 15752 31340 15804 31346
rect 15752 31282 15804 31288
rect 16028 31340 16080 31346
rect 16028 31282 16080 31288
rect 15396 30382 15516 30410
rect 15200 30252 15252 30258
rect 15200 30194 15252 30200
rect 15292 30184 15344 30190
rect 15292 30126 15344 30132
rect 15304 29782 15332 30126
rect 15292 29776 15344 29782
rect 15292 29718 15344 29724
rect 15488 29646 15516 30382
rect 15658 29744 15714 29753
rect 15658 29679 15714 29688
rect 15672 29646 15700 29679
rect 15108 29640 15160 29646
rect 15108 29582 15160 29588
rect 15476 29640 15528 29646
rect 15476 29582 15528 29588
rect 15660 29640 15712 29646
rect 15660 29582 15712 29588
rect 15016 29572 15068 29578
rect 15016 29514 15068 29520
rect 15028 26994 15056 29514
rect 15120 29345 15148 29582
rect 15106 29336 15162 29345
rect 15106 29271 15162 29280
rect 15120 28994 15148 29271
rect 15120 28966 15332 28994
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 15016 26988 15068 26994
rect 15016 26930 15068 26936
rect 15108 26852 15160 26858
rect 15108 26794 15160 26800
rect 15120 26518 15148 26794
rect 14924 26512 14976 26518
rect 14924 26454 14976 26460
rect 15108 26512 15160 26518
rect 15108 26454 15160 26460
rect 15108 25764 15160 25770
rect 15108 25706 15160 25712
rect 15120 25430 15148 25706
rect 15212 25430 15240 28018
rect 15304 26382 15332 28966
rect 15488 27962 15516 29582
rect 15396 27934 15516 27962
rect 15764 27946 15792 31282
rect 15936 30592 15988 30598
rect 15936 30534 15988 30540
rect 15844 30116 15896 30122
rect 15844 30058 15896 30064
rect 15856 29646 15884 30058
rect 15844 29640 15896 29646
rect 15844 29582 15896 29588
rect 15844 28144 15896 28150
rect 15844 28086 15896 28092
rect 15752 27940 15804 27946
rect 15396 26994 15424 27934
rect 15752 27882 15804 27888
rect 15476 27872 15528 27878
rect 15476 27814 15528 27820
rect 15488 27062 15516 27814
rect 15568 27464 15620 27470
rect 15620 27412 15792 27418
rect 15568 27406 15792 27412
rect 15580 27390 15792 27406
rect 15568 27328 15620 27334
rect 15568 27270 15620 27276
rect 15476 27056 15528 27062
rect 15476 26998 15528 27004
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 15108 25424 15160 25430
rect 15108 25366 15160 25372
rect 15200 25424 15252 25430
rect 15200 25366 15252 25372
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 15200 24948 15252 24954
rect 15200 24890 15252 24896
rect 15212 24857 15240 24890
rect 15198 24848 15254 24857
rect 15198 24783 15254 24792
rect 14740 24744 14792 24750
rect 14924 24744 14976 24750
rect 14740 24686 14792 24692
rect 14844 24704 14924 24732
rect 14752 24342 14780 24686
rect 14740 24336 14792 24342
rect 14740 24278 14792 24284
rect 14844 23866 14872 24704
rect 14924 24686 14976 24692
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15120 24206 15148 24550
rect 15212 24342 15240 24783
rect 15200 24336 15252 24342
rect 15200 24278 15252 24284
rect 15304 24274 15332 26318
rect 15396 26296 15424 26930
rect 15476 26920 15528 26926
rect 15476 26862 15528 26868
rect 15488 26450 15516 26862
rect 15580 26790 15608 27270
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15580 26518 15608 26726
rect 15568 26512 15620 26518
rect 15568 26454 15620 26460
rect 15476 26444 15528 26450
rect 15476 26386 15528 26392
rect 15476 26308 15528 26314
rect 15396 26268 15476 26296
rect 15528 26268 15608 26296
rect 15476 26250 15528 26256
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15396 24410 15424 24754
rect 15384 24404 15436 24410
rect 15384 24346 15436 24352
rect 15580 24342 15608 26268
rect 15672 25294 15700 26930
rect 15764 26382 15792 27390
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 15568 24336 15620 24342
rect 15568 24278 15620 24284
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 14936 23730 14964 24142
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 15028 23798 15056 24074
rect 15016 23792 15068 23798
rect 15016 23734 15068 23740
rect 14924 23724 14976 23730
rect 14924 23666 14976 23672
rect 14832 23520 14884 23526
rect 14832 23462 14884 23468
rect 14648 23044 14700 23050
rect 14648 22986 14700 22992
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14188 22374 14240 22380
rect 14200 22030 14228 22374
rect 14384 22358 14596 22386
rect 14384 22098 14412 22358
rect 14372 22092 14424 22098
rect 14372 22034 14424 22040
rect 14188 22024 14240 22030
rect 14188 21966 14240 21972
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 14004 21616 14056 21622
rect 14004 21558 14056 21564
rect 14016 21078 14044 21558
rect 14200 21554 14228 21966
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14188 21548 14240 21554
rect 14372 21548 14424 21554
rect 14240 21508 14320 21536
rect 14188 21490 14240 21496
rect 14004 21072 14056 21078
rect 14004 21014 14056 21020
rect 13912 20936 13964 20942
rect 13912 20878 13964 20884
rect 13924 19310 13952 20878
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 14016 20534 14044 20810
rect 14108 20806 14136 21490
rect 14186 21040 14242 21049
rect 14186 20975 14242 20984
rect 14200 20942 14228 20975
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 14016 20058 14044 20470
rect 14108 20058 14136 20742
rect 14292 20602 14320 21508
rect 14372 21490 14424 21496
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 14016 19718 14044 19790
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13924 18426 13952 18838
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14016 18290 14044 19654
rect 14292 19378 14320 20538
rect 14384 19990 14412 21490
rect 14568 20806 14596 21898
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14660 20618 14688 22578
rect 14738 21720 14794 21729
rect 14738 21655 14740 21664
rect 14792 21655 14794 21664
rect 14740 21626 14792 21632
rect 14752 21146 14780 21626
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14568 20590 14688 20618
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14200 18426 14228 18566
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 15026 13860 16390
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13740 13258 13768 14962
rect 13832 14550 13860 14962
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13832 14074 13860 14486
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13648 12986 13676 13126
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13740 10062 13768 13194
rect 13832 13190 13860 13466
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12986 13860 13126
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13924 10266 13952 18158
rect 14200 17678 14228 18226
rect 14292 18086 14320 19314
rect 14568 19292 14596 20590
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14660 19553 14688 20470
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14646 19544 14702 19553
rect 14646 19479 14702 19488
rect 14476 19264 14596 19292
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 14016 17338 14044 17478
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14292 16794 14320 18022
rect 14476 17678 14504 19264
rect 14660 19242 14688 19479
rect 14752 19378 14780 19858
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14648 19236 14700 19242
rect 14648 19178 14700 19184
rect 14752 19122 14780 19314
rect 14568 19094 14780 19122
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14372 17604 14424 17610
rect 14372 17546 14424 17552
rect 14384 17066 14412 17546
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14200 15706 14228 16050
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14108 14618 14136 14962
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13740 9586 13768 9998
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13740 8294 13768 8978
rect 13832 8974 13860 9522
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13728 8288 13780 8294
rect 13648 8248 13728 8276
rect 13648 7954 13676 8248
rect 13728 8230 13780 8236
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13544 7268 13596 7274
rect 13544 7210 13596 7216
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12912 6798 12940 7142
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12452 6310 12572 6338
rect 12360 6186 12480 6202
rect 12348 6180 12480 6186
rect 12400 6174 12480 6180
rect 12348 6122 12400 6128
rect 12452 5710 12480 6174
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11716 5302 11744 5510
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11164 4826 11192 4966
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 12176 4690 12204 5306
rect 12544 5302 12572 6310
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12636 5710 12664 6190
rect 13556 5846 13584 7210
rect 13648 7002 13676 7754
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13648 6322 13676 6938
rect 13740 6866 13768 8026
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12544 5030 12572 5238
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 12544 4554 12572 4966
rect 12636 4826 12664 5646
rect 12992 5636 13044 5642
rect 12992 5578 13044 5584
rect 13004 5166 13032 5578
rect 13832 5574 13860 6598
rect 13924 6458 13952 9318
rect 14016 7954 14044 14214
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 10742 14136 10950
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14108 9178 14136 9522
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 14200 5914 14228 15642
rect 14292 15008 14320 16730
rect 14384 15502 14412 17002
rect 14476 16250 14504 17614
rect 14568 17134 14596 19094
rect 14738 18320 14794 18329
rect 14738 18255 14794 18264
rect 14752 18222 14780 18255
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14660 17746 14688 18022
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14568 16590 14596 17070
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14568 16250 14596 16526
rect 14464 16244 14516 16250
rect 14464 16186 14516 16192
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14568 16114 14596 16186
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14568 15162 14596 16050
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14372 15020 14424 15026
rect 14292 14980 14372 15008
rect 14372 14962 14424 14968
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14292 14278 14320 14826
rect 14384 14521 14412 14962
rect 14660 14958 14688 15438
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14370 14512 14426 14521
rect 14370 14447 14372 14456
rect 14424 14447 14426 14456
rect 14372 14418 14424 14424
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 11694 14320 14214
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14660 13258 14688 13874
rect 14752 13530 14780 17818
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14844 12730 14872 23462
rect 14936 21690 14964 23666
rect 15028 23474 15056 23734
rect 15120 23730 15148 24142
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15488 23730 15516 24006
rect 15672 23866 15700 25230
rect 15752 24880 15804 24886
rect 15752 24822 15804 24828
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15108 23724 15160 23730
rect 15108 23666 15160 23672
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15028 23446 15240 23474
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 15028 23118 15056 23258
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15120 21962 15148 23054
rect 15212 22778 15240 23446
rect 15304 23322 15332 23666
rect 15292 23316 15344 23322
rect 15292 23258 15344 23264
rect 15568 23180 15620 23186
rect 15568 23122 15620 23128
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15200 22772 15252 22778
rect 15396 22760 15424 23054
rect 15580 22982 15608 23122
rect 15568 22976 15620 22982
rect 15568 22918 15620 22924
rect 15200 22714 15252 22720
rect 15304 22732 15424 22760
rect 15476 22772 15528 22778
rect 15304 22114 15332 22732
rect 15476 22714 15528 22720
rect 15384 22160 15436 22166
rect 15304 22108 15384 22114
rect 15304 22102 15436 22108
rect 15304 22086 15424 22102
rect 15108 21956 15160 21962
rect 15108 21898 15160 21904
rect 15198 21720 15254 21729
rect 14924 21684 14976 21690
rect 15198 21655 15254 21664
rect 14924 21626 14976 21632
rect 15212 21554 15240 21655
rect 15304 21554 15332 22086
rect 15488 22030 15516 22714
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15580 22030 15608 22578
rect 15672 22098 15700 23122
rect 15660 22092 15712 22098
rect 15660 22034 15712 22040
rect 15384 22024 15436 22030
rect 15384 21966 15436 21972
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15568 22024 15620 22030
rect 15764 22012 15792 24822
rect 15856 24410 15884 28086
rect 15948 26489 15976 30534
rect 16040 29578 16068 31282
rect 16132 30818 16160 31350
rect 16212 31340 16264 31346
rect 16212 31282 16264 31288
rect 16224 31210 16252 31282
rect 16316 31249 16344 33934
rect 16396 33856 16448 33862
rect 16396 33798 16448 33804
rect 16408 32910 16436 33798
rect 16500 33590 16528 33952
rect 16488 33584 16540 33590
rect 16488 33526 16540 33532
rect 16396 32904 16448 32910
rect 16396 32846 16448 32852
rect 16408 32502 16436 32846
rect 16396 32496 16448 32502
rect 16396 32438 16448 32444
rect 16408 31822 16436 32438
rect 16396 31816 16448 31822
rect 16396 31758 16448 31764
rect 16396 31408 16448 31414
rect 16592 31396 16620 37828
rect 16856 37810 16908 37816
rect 17224 37868 17276 37874
rect 17224 37810 17276 37816
rect 17684 37868 17736 37874
rect 17684 37810 17736 37816
rect 17868 37868 17920 37874
rect 17868 37810 17920 37816
rect 20364 37862 20668 37890
rect 20824 37874 20852 38286
rect 20996 38208 21048 38214
rect 20996 38150 21048 38156
rect 21008 38010 21036 38150
rect 21284 38010 21312 38286
rect 22008 38208 22060 38214
rect 22008 38150 22060 38156
rect 24032 38208 24084 38214
rect 24032 38150 24084 38156
rect 20996 38004 21048 38010
rect 20996 37946 21048 37952
rect 21272 38004 21324 38010
rect 21272 37946 21324 37952
rect 16764 36372 16816 36378
rect 16764 36314 16816 36320
rect 16776 36174 16804 36314
rect 16868 36174 16896 37810
rect 17132 37120 17184 37126
rect 17132 37062 17184 37068
rect 17040 36712 17092 36718
rect 17040 36654 17092 36660
rect 16672 36168 16724 36174
rect 16672 36110 16724 36116
rect 16764 36168 16816 36174
rect 16764 36110 16816 36116
rect 16856 36168 16908 36174
rect 16856 36110 16908 36116
rect 16684 33658 16712 36110
rect 17052 36106 17080 36654
rect 17144 36310 17172 37062
rect 17132 36304 17184 36310
rect 17132 36246 17184 36252
rect 17144 36106 17172 36246
rect 17236 36174 17264 37810
rect 17500 36780 17552 36786
rect 17500 36722 17552 36728
rect 17224 36168 17276 36174
rect 17224 36110 17276 36116
rect 17040 36100 17092 36106
rect 17040 36042 17092 36048
rect 17132 36100 17184 36106
rect 17132 36042 17184 36048
rect 16764 34672 16816 34678
rect 16764 34614 16816 34620
rect 16776 33946 16804 34614
rect 17132 34604 17184 34610
rect 17132 34546 17184 34552
rect 16856 34400 16908 34406
rect 16856 34342 16908 34348
rect 16948 34400 17000 34406
rect 16948 34342 17000 34348
rect 17040 34400 17092 34406
rect 17040 34342 17092 34348
rect 16868 34202 16896 34342
rect 16960 34202 16988 34342
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 16948 34196 17000 34202
rect 16948 34138 17000 34144
rect 16856 34060 16908 34066
rect 17052 34048 17080 34342
rect 17144 34202 17172 34546
rect 17132 34196 17184 34202
rect 17132 34138 17184 34144
rect 16908 34020 17080 34048
rect 16856 34002 16908 34008
rect 17132 33992 17184 33998
rect 16776 33918 16896 33946
rect 16672 33652 16724 33658
rect 16672 33594 16724 33600
rect 16684 32774 16712 33594
rect 16672 32768 16724 32774
rect 16672 32710 16724 32716
rect 16764 32224 16816 32230
rect 16764 32166 16816 32172
rect 16672 31476 16724 31482
rect 16672 31418 16724 31424
rect 16448 31368 16620 31396
rect 16396 31350 16448 31356
rect 16302 31240 16358 31249
rect 16212 31204 16264 31210
rect 16302 31175 16358 31184
rect 16212 31146 16264 31152
rect 16224 30938 16252 31146
rect 16212 30932 16264 30938
rect 16212 30874 16264 30880
rect 16132 30790 16252 30818
rect 16120 30252 16172 30258
rect 16120 30194 16172 30200
rect 16132 29646 16160 30194
rect 16120 29640 16172 29646
rect 16120 29582 16172 29588
rect 16028 29572 16080 29578
rect 16028 29514 16080 29520
rect 16040 29102 16068 29514
rect 16028 29096 16080 29102
rect 16028 29038 16080 29044
rect 16224 28558 16252 30790
rect 16316 30598 16344 31175
rect 16304 30592 16356 30598
rect 16304 30534 16356 30540
rect 16408 30297 16436 31350
rect 16684 31210 16712 31418
rect 16672 31204 16724 31210
rect 16672 31146 16724 31152
rect 16488 31136 16540 31142
rect 16488 31078 16540 31084
rect 16394 30288 16450 30297
rect 16500 30258 16528 31078
rect 16684 30734 16712 31146
rect 16580 30728 16632 30734
rect 16580 30670 16632 30676
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16394 30223 16450 30232
rect 16488 30252 16540 30258
rect 16408 30138 16436 30223
rect 16488 30194 16540 30200
rect 16408 30110 16528 30138
rect 16396 29572 16448 29578
rect 16396 29514 16448 29520
rect 16304 28688 16356 28694
rect 16304 28630 16356 28636
rect 16120 28552 16172 28558
rect 16120 28494 16172 28500
rect 16212 28552 16264 28558
rect 16212 28494 16264 28500
rect 16132 28218 16160 28494
rect 16120 28212 16172 28218
rect 16120 28154 16172 28160
rect 16028 28076 16080 28082
rect 16028 28018 16080 28024
rect 16040 27674 16068 28018
rect 16120 27872 16172 27878
rect 16120 27814 16172 27820
rect 16028 27668 16080 27674
rect 16028 27610 16080 27616
rect 16132 27470 16160 27814
rect 16120 27464 16172 27470
rect 16120 27406 16172 27412
rect 15934 26480 15990 26489
rect 15934 26415 15990 26424
rect 15948 26314 15976 26415
rect 15936 26308 15988 26314
rect 15936 26250 15988 26256
rect 15844 24404 15896 24410
rect 15844 24346 15896 24352
rect 15856 24206 15884 24346
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15948 23866 15976 26250
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 16040 23662 16068 24142
rect 16028 23656 16080 23662
rect 16028 23598 16080 23604
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15856 22778 15884 23054
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 16040 22506 16068 23258
rect 16132 23186 16160 27406
rect 16316 27130 16344 28630
rect 16304 27124 16356 27130
rect 16304 27066 16356 27072
rect 16212 25288 16264 25294
rect 16212 25230 16264 25236
rect 16224 23526 16252 25230
rect 16316 24886 16344 27066
rect 16408 26994 16436 29514
rect 16500 28558 16528 30110
rect 16592 29850 16620 30670
rect 16672 30592 16724 30598
rect 16776 30580 16804 32166
rect 16868 31385 16896 33918
rect 17052 33940 17132 33946
rect 17052 33934 17184 33940
rect 17052 33918 17172 33934
rect 16948 33856 17000 33862
rect 17052 33844 17080 33918
rect 17000 33816 17080 33844
rect 16948 33798 17000 33804
rect 17052 32502 17080 33816
rect 17137 33856 17189 33862
rect 17137 33798 17189 33804
rect 17040 32496 17092 32502
rect 17040 32438 17092 32444
rect 16854 31376 16910 31385
rect 16854 31311 16910 31320
rect 16868 30870 16896 31311
rect 16856 30864 16908 30870
rect 16856 30806 16908 30812
rect 16868 30734 16896 30806
rect 16948 30796 17000 30802
rect 16948 30738 17000 30744
rect 16856 30728 16908 30734
rect 16856 30670 16908 30676
rect 16776 30552 16896 30580
rect 16672 30534 16724 30540
rect 16684 30190 16712 30534
rect 16672 30184 16724 30190
rect 16672 30126 16724 30132
rect 16764 30184 16816 30190
rect 16764 30126 16816 30132
rect 16776 30036 16804 30126
rect 16684 30008 16804 30036
rect 16868 30036 16896 30552
rect 16960 30190 16988 30738
rect 16948 30184 17000 30190
rect 16948 30126 17000 30132
rect 16868 30008 16988 30036
rect 16580 29844 16632 29850
rect 16580 29786 16632 29792
rect 16684 29170 16712 30008
rect 16960 29510 16988 30008
rect 17052 29510 17080 32438
rect 17144 32230 17172 33798
rect 17236 32910 17264 36110
rect 17408 36032 17460 36038
rect 17406 36000 17408 36009
rect 17460 36000 17462 36009
rect 17406 35935 17462 35944
rect 17512 35850 17540 36722
rect 17592 36100 17644 36106
rect 17592 36042 17644 36048
rect 17420 35822 17540 35850
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 17328 34746 17356 35022
rect 17316 34740 17368 34746
rect 17316 34682 17368 34688
rect 17316 34196 17368 34202
rect 17316 34138 17368 34144
rect 17328 33998 17356 34138
rect 17420 34082 17448 35822
rect 17604 34746 17632 36042
rect 17592 34740 17644 34746
rect 17592 34682 17644 34688
rect 17696 34082 17724 37810
rect 17880 37466 17908 37810
rect 19984 37800 20036 37806
rect 19154 37768 19210 37777
rect 20364 37754 20392 37862
rect 20036 37748 20392 37754
rect 19984 37742 20392 37748
rect 20444 37800 20496 37806
rect 20444 37742 20496 37748
rect 19294 37732 19346 37738
rect 19210 37712 19294 37720
rect 19154 37703 19294 37712
rect 19168 37692 19294 37703
rect 19996 37726 20392 37742
rect 19294 37674 19346 37680
rect 17960 37664 18012 37670
rect 17960 37606 18012 37612
rect 17868 37460 17920 37466
rect 17868 37402 17920 37408
rect 17972 37346 18000 37606
rect 17880 37330 18000 37346
rect 17868 37324 18000 37330
rect 17920 37318 18000 37324
rect 17868 37266 17920 37272
rect 18420 37256 18472 37262
rect 18420 37198 18472 37204
rect 17776 37188 17828 37194
rect 17776 37130 17828 37136
rect 17788 36378 17816 37130
rect 18432 36786 18460 37198
rect 18512 37120 18564 37126
rect 18512 37062 18564 37068
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 17960 36576 18012 36582
rect 17960 36518 18012 36524
rect 17776 36372 17828 36378
rect 17776 36314 17828 36320
rect 17972 36242 18000 36518
rect 17960 36236 18012 36242
rect 17960 36178 18012 36184
rect 17868 36168 17920 36174
rect 17868 36110 17920 36116
rect 18052 36168 18104 36174
rect 18052 36110 18104 36116
rect 17420 34054 17540 34082
rect 17316 33992 17368 33998
rect 17316 33934 17368 33940
rect 17316 33856 17368 33862
rect 17316 33798 17368 33804
rect 17328 33658 17356 33798
rect 17316 33652 17368 33658
rect 17316 33594 17368 33600
rect 17328 33114 17356 33594
rect 17512 33402 17540 34054
rect 17604 34054 17724 34082
rect 17776 34128 17828 34134
rect 17776 34070 17828 34076
rect 17604 33538 17632 34054
rect 17684 33992 17736 33998
rect 17684 33934 17736 33940
rect 17696 33658 17724 33934
rect 17684 33652 17736 33658
rect 17684 33594 17736 33600
rect 17604 33510 17724 33538
rect 17788 33522 17816 34070
rect 17420 33374 17540 33402
rect 17592 33380 17644 33386
rect 17316 33108 17368 33114
rect 17316 33050 17368 33056
rect 17224 32904 17276 32910
rect 17224 32846 17276 32852
rect 17132 32224 17184 32230
rect 17132 32166 17184 32172
rect 17236 31754 17264 32846
rect 17224 31748 17276 31754
rect 17224 31690 17276 31696
rect 17236 31210 17264 31690
rect 17328 31346 17356 33050
rect 17316 31340 17368 31346
rect 17316 31282 17368 31288
rect 17224 31204 17276 31210
rect 17224 31146 17276 31152
rect 17132 30864 17184 30870
rect 17132 30806 17184 30812
rect 16764 29504 16816 29510
rect 16764 29446 16816 29452
rect 16856 29504 16908 29510
rect 16856 29446 16908 29452
rect 16948 29504 17000 29510
rect 16948 29446 17000 29452
rect 17040 29504 17092 29510
rect 17040 29446 17092 29452
rect 16776 29306 16804 29446
rect 16764 29300 16816 29306
rect 16764 29242 16816 29248
rect 16868 29170 16896 29446
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16488 28552 16540 28558
rect 16488 28494 16540 28500
rect 16856 28484 16908 28490
rect 16856 28426 16908 28432
rect 16488 28416 16540 28422
rect 16488 28358 16540 28364
rect 16500 27305 16528 28358
rect 16580 28212 16632 28218
rect 16580 28154 16632 28160
rect 16592 27470 16620 28154
rect 16868 28150 16896 28426
rect 16856 28144 16908 28150
rect 16856 28086 16908 28092
rect 16764 28076 16816 28082
rect 16764 28018 16816 28024
rect 16776 27470 16804 28018
rect 16854 27568 16910 27577
rect 16854 27503 16910 27512
rect 16580 27464 16632 27470
rect 16580 27406 16632 27412
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16764 27464 16816 27470
rect 16764 27406 16816 27412
rect 16486 27296 16542 27305
rect 16486 27231 16542 27240
rect 16684 27130 16712 27406
rect 16868 27334 16896 27503
rect 16856 27328 16908 27334
rect 16856 27270 16908 27276
rect 16960 27130 16988 29446
rect 16672 27124 16724 27130
rect 16672 27066 16724 27072
rect 16948 27124 17000 27130
rect 16948 27066 17000 27072
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 16486 26344 16542 26353
rect 16408 26302 16486 26330
rect 16304 24880 16356 24886
rect 16304 24822 16356 24828
rect 16408 24154 16436 26302
rect 16486 26279 16542 26288
rect 16776 25974 16804 26930
rect 16960 26926 16988 27066
rect 17052 26994 17080 29446
rect 17144 27606 17172 30806
rect 17224 30592 17276 30598
rect 17224 30534 17276 30540
rect 17236 30190 17264 30534
rect 17224 30184 17276 30190
rect 17224 30126 17276 30132
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17132 27600 17184 27606
rect 17132 27542 17184 27548
rect 17236 27452 17264 29106
rect 17328 28082 17356 31282
rect 17420 30734 17448 33374
rect 17592 33322 17644 33328
rect 17500 32496 17552 32502
rect 17604 32484 17632 33322
rect 17696 33153 17724 33510
rect 17776 33516 17828 33522
rect 17776 33458 17828 33464
rect 17682 33144 17738 33153
rect 17682 33079 17738 33088
rect 17696 32570 17724 33079
rect 17684 32564 17736 32570
rect 17684 32506 17736 32512
rect 17552 32456 17632 32484
rect 17500 32438 17552 32444
rect 17408 30728 17460 30734
rect 17408 30670 17460 30676
rect 17408 30048 17460 30054
rect 17408 29990 17460 29996
rect 17420 29850 17448 29990
rect 17408 29844 17460 29850
rect 17408 29786 17460 29792
rect 17512 29170 17540 32438
rect 17592 32292 17644 32298
rect 17592 32234 17644 32240
rect 17604 32026 17632 32234
rect 17592 32020 17644 32026
rect 17592 31962 17644 31968
rect 17880 31634 17908 36110
rect 17960 35624 18012 35630
rect 17960 35566 18012 35572
rect 17972 34513 18000 35566
rect 17958 34504 18014 34513
rect 17958 34439 18014 34448
rect 18064 34406 18092 36110
rect 18144 35012 18196 35018
rect 18144 34954 18196 34960
rect 18052 34400 18104 34406
rect 18052 34342 18104 34348
rect 17960 34196 18012 34202
rect 17960 34138 18012 34144
rect 17972 34105 18000 34138
rect 17958 34096 18014 34105
rect 17958 34031 18014 34040
rect 18064 33930 18092 34342
rect 17960 33924 18012 33930
rect 17960 33866 18012 33872
rect 18052 33924 18104 33930
rect 18052 33866 18104 33872
rect 17972 33810 18000 33866
rect 18156 33810 18184 34954
rect 18420 33992 18472 33998
rect 18420 33934 18472 33940
rect 18236 33924 18288 33930
rect 18236 33866 18288 33872
rect 17972 33782 18184 33810
rect 18156 33386 18184 33782
rect 18144 33380 18196 33386
rect 18064 33340 18144 33368
rect 17958 31920 18014 31929
rect 17958 31855 17960 31864
rect 18012 31855 18014 31864
rect 17960 31826 18012 31832
rect 17788 31606 17908 31634
rect 17788 31346 17816 31606
rect 17866 31512 17922 31521
rect 17866 31447 17922 31456
rect 17880 31414 17908 31447
rect 17868 31408 17920 31414
rect 17868 31350 17920 31356
rect 18064 31346 18092 33340
rect 18144 33322 18196 33328
rect 18248 32842 18276 33866
rect 18328 33856 18380 33862
rect 18328 33798 18380 33804
rect 18340 33114 18368 33798
rect 18432 33318 18460 33934
rect 18420 33312 18472 33318
rect 18420 33254 18472 33260
rect 18328 33108 18380 33114
rect 18328 33050 18380 33056
rect 18236 32836 18288 32842
rect 18236 32778 18288 32784
rect 18420 32428 18472 32434
rect 18420 32370 18472 32376
rect 18432 32065 18460 32370
rect 18418 32056 18474 32065
rect 18144 32020 18196 32026
rect 18418 31991 18474 32000
rect 18144 31962 18196 31968
rect 18156 31754 18184 31962
rect 18328 31884 18380 31890
rect 18328 31826 18380 31832
rect 18156 31726 18276 31754
rect 18144 31680 18196 31686
rect 18144 31622 18196 31628
rect 17592 31340 17644 31346
rect 17592 31282 17644 31288
rect 17684 31340 17736 31346
rect 17684 31282 17736 31288
rect 17776 31340 17828 31346
rect 17776 31282 17828 31288
rect 18052 31340 18104 31346
rect 18052 31282 18104 31288
rect 17604 30938 17632 31282
rect 17592 30932 17644 30938
rect 17592 30874 17644 30880
rect 17592 30728 17644 30734
rect 17592 30670 17644 30676
rect 17500 29164 17552 29170
rect 17500 29106 17552 29112
rect 17316 28076 17368 28082
rect 17316 28018 17368 28024
rect 17316 27872 17368 27878
rect 17316 27814 17368 27820
rect 17408 27872 17460 27878
rect 17408 27814 17460 27820
rect 17144 27424 17264 27452
rect 17040 26988 17092 26994
rect 17040 26930 17092 26936
rect 16948 26920 17000 26926
rect 16948 26862 17000 26868
rect 17144 26858 17172 27424
rect 17328 27316 17356 27814
rect 17420 27470 17448 27814
rect 17604 27606 17632 30670
rect 17696 29753 17724 31282
rect 17682 29744 17738 29753
rect 17682 29679 17738 29688
rect 17684 29164 17736 29170
rect 17684 29106 17736 29112
rect 17696 28937 17724 29106
rect 17682 28928 17738 28937
rect 17682 28863 17738 28872
rect 17696 27878 17724 28863
rect 17684 27872 17736 27878
rect 17684 27814 17736 27820
rect 17592 27600 17644 27606
rect 17592 27542 17644 27548
rect 17684 27600 17736 27606
rect 17684 27542 17736 27548
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17500 27464 17552 27470
rect 17500 27406 17552 27412
rect 17512 27316 17540 27406
rect 17328 27288 17540 27316
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17132 26852 17184 26858
rect 17132 26794 17184 26800
rect 16948 26784 17000 26790
rect 16948 26726 17000 26732
rect 16960 26382 16988 26726
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 16764 25968 16816 25974
rect 16764 25910 16816 25916
rect 16580 25832 16632 25838
rect 16580 25774 16632 25780
rect 16408 24126 16528 24154
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 16120 23180 16172 23186
rect 16120 23122 16172 23128
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 16028 22500 16080 22506
rect 16028 22442 16080 22448
rect 16132 22030 16160 22646
rect 16120 22024 16172 22030
rect 15764 21984 15884 22012
rect 15568 21966 15620 21972
rect 15396 21554 15424 21966
rect 15200 21548 15252 21554
rect 15120 21508 15200 21536
rect 14924 20868 14976 20874
rect 14924 20810 14976 20816
rect 14936 15706 14964 20810
rect 15120 20534 15148 21508
rect 15200 21490 15252 21496
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 15120 17746 15148 20334
rect 15212 17882 15240 20742
rect 15396 18426 15424 21490
rect 15488 21146 15516 21966
rect 15476 21140 15528 21146
rect 15476 21082 15528 21088
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15488 19854 15516 20742
rect 15580 20602 15608 21966
rect 15856 21876 15884 21984
rect 16120 21966 16172 21972
rect 15856 21848 16068 21876
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15672 20602 15700 20742
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15488 18630 15516 19790
rect 15580 19334 15608 20402
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15672 19514 15700 19790
rect 15856 19514 15884 19926
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 15580 19306 15700 19334
rect 15672 18737 15700 19306
rect 15658 18728 15714 18737
rect 15658 18663 15714 18672
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15488 18154 15516 18566
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15120 15978 15148 17682
rect 15396 17610 15424 18022
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15396 16590 15424 17546
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15108 15972 15160 15978
rect 15108 15914 15160 15920
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14936 12850 14964 15098
rect 15120 15042 15148 15914
rect 15028 15014 15148 15042
rect 15488 15026 15516 18090
rect 15580 17338 15608 18158
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15580 17202 15608 17274
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15672 16658 15700 18663
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15764 17746 15792 18566
rect 15948 18222 15976 21558
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15752 17604 15804 17610
rect 15752 17546 15804 17552
rect 15764 17134 15792 17546
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15660 16652 15712 16658
rect 15580 16612 15660 16640
rect 15580 16454 15608 16612
rect 15660 16594 15712 16600
rect 15856 16590 15884 17614
rect 15844 16584 15896 16590
rect 15764 16544 15844 16572
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15476 15020 15528 15026
rect 15028 14958 15056 15014
rect 15476 14962 15528 14968
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 15028 14482 15056 14894
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15212 13258 15240 13874
rect 15304 13530 15332 14350
rect 15580 13734 15608 15642
rect 15764 15570 15792 16544
rect 15844 16526 15896 16532
rect 15844 15700 15896 15706
rect 15948 15688 15976 18158
rect 15896 15660 15976 15688
rect 15844 15642 15896 15648
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 15936 15496 15988 15502
rect 15856 15456 15936 15484
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15764 14278 15792 15370
rect 15856 14618 15884 15456
rect 15936 15438 15988 15444
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15948 14278 15976 14962
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15212 12986 15240 13194
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14844 12702 15240 12730
rect 15108 12640 15160 12646
rect 15028 12588 15108 12594
rect 15028 12582 15160 12588
rect 15028 12566 15148 12582
rect 15028 12434 15056 12566
rect 15212 12458 15240 12702
rect 14752 12406 15056 12434
rect 15120 12430 15240 12458
rect 14752 12238 14780 12406
rect 15120 12322 15148 12430
rect 15028 12294 15148 12322
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14476 11354 14504 11834
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14844 11218 14872 11698
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 15028 10690 15056 12294
rect 15304 12186 15332 13126
rect 15476 12844 15528 12850
rect 15212 12158 15332 12186
rect 15396 12804 15476 12832
rect 15028 10662 15148 10690
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14384 9654 14412 10202
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14384 8974 14412 9590
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14660 8634 14688 8774
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14292 5642 14320 7278
rect 14660 6390 14688 7414
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 13648 5302 13676 5510
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 14384 4146 14412 5510
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14476 4282 14504 4490
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 12530 4040 12586 4049
rect 12530 3975 12586 3984
rect 13174 4040 13230 4049
rect 13174 3975 13230 3984
rect 12544 3058 12572 3975
rect 13188 3058 13216 3975
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 13004 2446 13032 2790
rect 14752 2774 14780 8774
rect 14936 8537 14964 8774
rect 14922 8528 14978 8537
rect 14922 8463 14978 8472
rect 15028 8430 15056 8910
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14936 5778 14964 7142
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 15120 3058 15148 10662
rect 15212 10656 15240 12158
rect 15292 12096 15344 12102
rect 15396 12084 15424 12804
rect 15476 12786 15528 12792
rect 15580 12434 15608 13126
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15344 12056 15424 12084
rect 15292 12038 15344 12044
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15304 11286 15332 11630
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 15292 10668 15344 10674
rect 15212 10628 15292 10656
rect 15292 10610 15344 10616
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15212 9024 15240 9454
rect 15304 9178 15332 9590
rect 15396 9586 15424 12056
rect 15488 12406 15608 12434
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15384 9036 15436 9042
rect 15212 8996 15384 9024
rect 15384 8978 15436 8984
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15396 7546 15424 7686
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15212 6118 15240 6734
rect 15304 6322 15332 7346
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15396 6322 15424 7278
rect 15488 7206 15516 12406
rect 15672 11914 15700 12718
rect 15580 11886 15700 11914
rect 15580 11694 15608 11886
rect 15660 11824 15712 11830
rect 15660 11766 15712 11772
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15580 11150 15608 11494
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15672 9518 15700 11766
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15764 10810 15792 11086
rect 15948 11014 15976 14214
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15672 8294 15700 9454
rect 15764 8974 15792 10746
rect 15948 10742 15976 10950
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 16040 9466 16068 21848
rect 16132 21729 16160 21966
rect 16224 21894 16252 23462
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 16316 22030 16344 22510
rect 16396 22160 16448 22166
rect 16396 22102 16448 22108
rect 16408 22030 16436 22102
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 16212 21888 16264 21894
rect 16212 21830 16264 21836
rect 16118 21720 16174 21729
rect 16118 21655 16174 21664
rect 16316 21622 16344 21966
rect 16304 21616 16356 21622
rect 16304 21558 16356 21564
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16132 20398 16160 20538
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 16132 20058 16160 20334
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16316 19854 16344 20198
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16224 19514 16252 19790
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16120 17672 16172 17678
rect 16224 17660 16252 19450
rect 16316 19446 16344 19790
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16172 17632 16252 17660
rect 16120 17614 16172 17620
rect 16132 15026 16160 17614
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16224 15026 16252 17274
rect 16316 16454 16344 19382
rect 16408 18290 16436 19790
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16316 14958 16344 16390
rect 16408 16250 16436 16390
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16408 15570 16436 16050
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16408 15162 16436 15506
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16408 14414 16436 14758
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16500 12866 16528 24126
rect 16592 22658 16620 25774
rect 17144 25430 17172 26794
rect 17132 25424 17184 25430
rect 17132 25366 17184 25372
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16776 24886 16804 25094
rect 16960 24954 16988 25230
rect 16948 24948 17000 24954
rect 16948 24890 17000 24896
rect 16764 24880 16816 24886
rect 16764 24822 16816 24828
rect 16776 24274 16804 24822
rect 16856 24676 16908 24682
rect 16856 24618 16908 24624
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16868 23798 16896 24618
rect 16948 24132 17000 24138
rect 17052 24120 17080 25230
rect 17132 25152 17184 25158
rect 17132 25094 17184 25100
rect 17144 24818 17172 25094
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 17144 24342 17172 24754
rect 17132 24336 17184 24342
rect 17132 24278 17184 24284
rect 17000 24092 17080 24120
rect 16948 24074 17000 24080
rect 17052 23866 17080 24092
rect 16948 23860 17000 23866
rect 16948 23802 17000 23808
rect 17040 23860 17092 23866
rect 17040 23802 17092 23808
rect 16856 23792 16908 23798
rect 16856 23734 16908 23740
rect 16764 23724 16816 23730
rect 16764 23666 16816 23672
rect 16776 22710 16804 23666
rect 16764 22704 16816 22710
rect 16592 22630 16712 22658
rect 16764 22646 16816 22652
rect 16580 21616 16632 21622
rect 16580 21558 16632 21564
rect 16592 21418 16620 21558
rect 16580 21412 16632 21418
rect 16580 21354 16632 21360
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16592 19786 16620 19926
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16592 16794 16620 17682
rect 16684 17082 16712 22630
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16764 22500 16816 22506
rect 16764 22442 16816 22448
rect 16776 22166 16804 22442
rect 16764 22160 16816 22166
rect 16764 22102 16816 22108
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16776 19242 16804 21966
rect 16868 20058 16896 22578
rect 16960 22166 16988 23802
rect 17236 23746 17264 26930
rect 17316 26852 17368 26858
rect 17316 26794 17368 26800
rect 17328 26586 17356 26794
rect 17500 26784 17552 26790
rect 17500 26726 17552 26732
rect 17316 26580 17368 26586
rect 17316 26522 17368 26528
rect 17512 26382 17540 26726
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17316 26240 17368 26246
rect 17314 26208 17316 26217
rect 17368 26208 17370 26217
rect 17314 26143 17370 26152
rect 17604 24954 17632 27542
rect 17696 27470 17724 27542
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 17788 27418 17816 31282
rect 17868 31136 17920 31142
rect 17868 31078 17920 31084
rect 17880 30054 17908 31078
rect 18052 30864 18104 30870
rect 18052 30806 18104 30812
rect 17960 30592 18012 30598
rect 17960 30534 18012 30540
rect 17868 30048 17920 30054
rect 17868 29990 17920 29996
rect 17972 29617 18000 30534
rect 18064 30394 18092 30806
rect 18156 30598 18184 31622
rect 18144 30592 18196 30598
rect 18144 30534 18196 30540
rect 18052 30388 18104 30394
rect 18052 30330 18104 30336
rect 18248 29730 18276 31726
rect 18340 31226 18368 31826
rect 18524 31754 18552 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19984 36780 20036 36786
rect 19984 36722 20036 36728
rect 19156 36712 19208 36718
rect 19156 36654 19208 36660
rect 19064 36100 19116 36106
rect 19064 36042 19116 36048
rect 18604 36032 18656 36038
rect 18604 35974 18656 35980
rect 18616 35766 18644 35974
rect 18604 35760 18656 35766
rect 18604 35702 18656 35708
rect 18880 35692 18932 35698
rect 18880 35634 18932 35640
rect 18696 35488 18748 35494
rect 18696 35430 18748 35436
rect 18602 33960 18658 33969
rect 18602 33895 18604 33904
rect 18656 33895 18658 33904
rect 18604 33866 18656 33872
rect 18708 33810 18736 35430
rect 18892 35290 18920 35634
rect 18880 35284 18932 35290
rect 18880 35226 18932 35232
rect 18788 35148 18840 35154
rect 18788 35090 18840 35096
rect 18800 33998 18828 35090
rect 18788 33992 18840 33998
rect 18788 33934 18840 33940
rect 19076 33930 19104 36042
rect 19168 34105 19196 36654
rect 19996 36310 20024 36722
rect 19984 36304 20036 36310
rect 19984 36246 20036 36252
rect 19340 36236 19392 36242
rect 19340 36178 19392 36184
rect 19352 35494 19380 36178
rect 19996 36106 20024 36246
rect 19984 36100 20036 36106
rect 19984 36042 20036 36048
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 20088 35816 20116 37726
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 20180 36009 20208 37198
rect 20456 36009 20484 37742
rect 20640 37720 20668 37862
rect 20812 37868 20864 37874
rect 20812 37810 20864 37816
rect 20720 37732 20772 37738
rect 20640 37692 20720 37720
rect 20720 37674 20772 37680
rect 20720 37188 20772 37194
rect 20720 37130 20772 37136
rect 20732 36922 20760 37130
rect 20720 36916 20772 36922
rect 20720 36858 20772 36864
rect 20720 36712 20772 36718
rect 20720 36654 20772 36660
rect 20536 36100 20588 36106
rect 20536 36042 20588 36048
rect 20166 36000 20222 36009
rect 20166 35935 20222 35944
rect 20442 36000 20498 36009
rect 20442 35935 20498 35944
rect 19904 35788 20116 35816
rect 19904 35737 19932 35788
rect 20444 35760 20496 35766
rect 19890 35728 19946 35737
rect 20444 35702 20496 35708
rect 19890 35663 19946 35672
rect 19984 35692 20036 35698
rect 19984 35634 20036 35640
rect 20076 35692 20128 35698
rect 20076 35634 20128 35640
rect 19340 35488 19392 35494
rect 19340 35430 19392 35436
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19246 34232 19302 34241
rect 19246 34167 19302 34176
rect 19154 34096 19210 34105
rect 19154 34031 19210 34040
rect 19064 33924 19116 33930
rect 19064 33866 19116 33872
rect 18616 33782 18736 33810
rect 18616 32434 18644 33782
rect 19064 33448 19116 33454
rect 19064 33390 19116 33396
rect 19076 33289 19104 33390
rect 19062 33280 19118 33289
rect 19062 33215 19118 33224
rect 18880 32972 18932 32978
rect 18880 32914 18932 32920
rect 18696 32904 18748 32910
rect 18696 32846 18748 32852
rect 18708 32434 18736 32846
rect 18604 32428 18656 32434
rect 18604 32370 18656 32376
rect 18696 32428 18748 32434
rect 18696 32370 18748 32376
rect 18708 32201 18736 32370
rect 18694 32192 18750 32201
rect 18694 32127 18750 32136
rect 18524 31726 18828 31754
rect 18696 31680 18748 31686
rect 18696 31622 18748 31628
rect 18708 31482 18736 31622
rect 18604 31476 18656 31482
rect 18604 31418 18656 31424
rect 18696 31476 18748 31482
rect 18696 31418 18748 31424
rect 18340 31198 18552 31226
rect 18328 31136 18380 31142
rect 18328 31078 18380 31084
rect 18340 30433 18368 31078
rect 18524 30666 18552 31198
rect 18512 30660 18564 30666
rect 18512 30602 18564 30608
rect 18326 30424 18382 30433
rect 18326 30359 18382 30368
rect 18524 30258 18552 30602
rect 18616 30258 18644 31418
rect 18800 31346 18828 31726
rect 18696 31340 18748 31346
rect 18696 31282 18748 31288
rect 18788 31340 18840 31346
rect 18788 31282 18840 31288
rect 18708 31226 18736 31282
rect 18892 31226 18920 32914
rect 19064 32836 19116 32842
rect 19064 32778 19116 32784
rect 19076 32434 19104 32778
rect 18972 32428 19024 32434
rect 18972 32370 19024 32376
rect 19064 32428 19116 32434
rect 19064 32370 19116 32376
rect 18984 32026 19012 32370
rect 18972 32020 19024 32026
rect 18972 31962 19024 31968
rect 19064 32020 19116 32026
rect 19064 31962 19116 31968
rect 19076 31754 19104 31962
rect 18708 31198 18920 31226
rect 18984 31726 19104 31754
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 18328 30184 18380 30190
rect 18380 30132 18460 30138
rect 18328 30126 18460 30132
rect 18340 30110 18460 30126
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 18340 29782 18368 29990
rect 18052 29708 18104 29714
rect 18052 29650 18104 29656
rect 18156 29702 18276 29730
rect 18328 29776 18380 29782
rect 18328 29718 18380 29724
rect 17958 29608 18014 29617
rect 17958 29543 18014 29552
rect 17972 29238 18000 29543
rect 17960 29232 18012 29238
rect 17960 29174 18012 29180
rect 18064 28937 18092 29650
rect 18156 29646 18184 29702
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 18050 28928 18106 28937
rect 18050 28863 18106 28872
rect 18050 28792 18106 28801
rect 18050 28727 18106 28736
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 17868 28484 17920 28490
rect 17868 28426 17920 28432
rect 17880 28082 17908 28426
rect 17868 28076 17920 28082
rect 17868 28018 17920 28024
rect 17866 27568 17922 27577
rect 17866 27503 17868 27512
rect 17920 27503 17922 27512
rect 17868 27474 17920 27480
rect 17788 27390 17908 27418
rect 17776 27328 17828 27334
rect 17682 27296 17738 27305
rect 17776 27270 17828 27276
rect 17682 27231 17738 27240
rect 17696 26994 17724 27231
rect 17788 26994 17816 27270
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17776 26988 17828 26994
rect 17776 26930 17828 26936
rect 17684 26784 17736 26790
rect 17684 26726 17736 26732
rect 17696 26586 17724 26726
rect 17684 26580 17736 26586
rect 17684 26522 17736 26528
rect 17880 26518 17908 27390
rect 17972 26518 18000 28494
rect 18064 27538 18092 28727
rect 18052 27532 18104 27538
rect 18052 27474 18104 27480
rect 18156 27470 18184 29582
rect 18432 29170 18460 30110
rect 18524 29730 18552 30194
rect 18708 30190 18736 31198
rect 18788 30592 18840 30598
rect 18788 30534 18840 30540
rect 18696 30184 18748 30190
rect 18696 30126 18748 30132
rect 18696 30048 18748 30054
rect 18696 29990 18748 29996
rect 18708 29782 18736 29990
rect 18696 29776 18748 29782
rect 18524 29702 18644 29730
rect 18696 29718 18748 29724
rect 18512 29640 18564 29646
rect 18512 29582 18564 29588
rect 18420 29164 18472 29170
rect 18420 29106 18472 29112
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 18328 28620 18380 28626
rect 18328 28562 18380 28568
rect 18236 27872 18288 27878
rect 18236 27814 18288 27820
rect 18144 27464 18196 27470
rect 18144 27406 18196 27412
rect 17868 26512 17920 26518
rect 17682 26480 17738 26489
rect 17868 26454 17920 26460
rect 17960 26512 18012 26518
rect 17960 26454 18012 26460
rect 17682 26415 17738 26424
rect 17776 26444 17828 26450
rect 17696 26314 17724 26415
rect 17776 26386 17828 26392
rect 17684 26308 17736 26314
rect 17684 26250 17736 26256
rect 17788 26217 17816 26386
rect 17774 26208 17830 26217
rect 17774 26143 17830 26152
rect 17776 25968 17828 25974
rect 17776 25910 17828 25916
rect 17788 25140 17816 25910
rect 17880 25430 17908 26454
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17868 25424 17920 25430
rect 17868 25366 17920 25372
rect 17868 25152 17920 25158
rect 17788 25112 17868 25140
rect 17868 25094 17920 25100
rect 17592 24948 17644 24954
rect 17592 24890 17644 24896
rect 17684 24880 17736 24886
rect 17684 24822 17736 24828
rect 17696 24750 17724 24822
rect 17880 24750 17908 25094
rect 17684 24744 17736 24750
rect 17684 24686 17736 24692
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17408 24676 17460 24682
rect 17408 24618 17460 24624
rect 17316 24336 17368 24342
rect 17316 24278 17368 24284
rect 17420 24290 17448 24618
rect 17696 24313 17724 24686
rect 17972 24682 18000 25842
rect 18156 25838 18184 27406
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18144 25696 18196 25702
rect 18144 25638 18196 25644
rect 18156 25362 18184 25638
rect 18248 25378 18276 27814
rect 18340 25906 18368 28562
rect 18432 28218 18460 28902
rect 18420 28212 18472 28218
rect 18420 28154 18472 28160
rect 18524 27554 18552 29582
rect 18616 29170 18644 29702
rect 18696 29640 18748 29646
rect 18696 29582 18748 29588
rect 18708 29306 18736 29582
rect 18696 29300 18748 29306
rect 18696 29242 18748 29248
rect 18604 29164 18656 29170
rect 18656 29124 18736 29152
rect 18604 29106 18656 29112
rect 18604 28960 18656 28966
rect 18604 28902 18656 28908
rect 18616 27690 18644 28902
rect 18708 27826 18736 29124
rect 18800 28218 18828 30534
rect 18984 30258 19012 31726
rect 19168 31346 19196 34031
rect 19260 33998 19288 34167
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19338 33824 19394 33833
rect 19338 33759 19394 33768
rect 19352 33658 19380 33759
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19340 33652 19392 33658
rect 19340 33594 19392 33600
rect 19708 33516 19760 33522
rect 19708 33458 19760 33464
rect 19616 33448 19668 33454
rect 19616 33390 19668 33396
rect 19432 33312 19484 33318
rect 19432 33254 19484 33260
rect 19444 32230 19472 33254
rect 19628 32978 19656 33390
rect 19616 32972 19668 32978
rect 19616 32914 19668 32920
rect 19720 32910 19748 33458
rect 19996 33386 20024 35634
rect 19892 33380 19944 33386
rect 19892 33322 19944 33328
rect 19984 33380 20036 33386
rect 19984 33322 20036 33328
rect 19708 32904 19760 32910
rect 19708 32846 19760 32852
rect 19904 32824 19932 33322
rect 19984 32836 20036 32842
rect 19904 32796 19984 32824
rect 19984 32778 20036 32784
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19432 32224 19484 32230
rect 19432 32166 19484 32172
rect 19984 32224 20036 32230
rect 19984 32166 20036 32172
rect 19156 31340 19208 31346
rect 19444 31328 19472 32166
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19996 31414 20024 32166
rect 19984 31408 20036 31414
rect 19984 31350 20036 31356
rect 19708 31340 19760 31346
rect 19444 31300 19708 31328
rect 19156 31282 19208 31288
rect 19708 31282 19760 31288
rect 19062 30832 19118 30841
rect 19062 30767 19118 30776
rect 19076 30734 19104 30767
rect 19064 30728 19116 30734
rect 19064 30670 19116 30676
rect 18972 30252 19024 30258
rect 18972 30194 19024 30200
rect 19064 30252 19116 30258
rect 19064 30194 19116 30200
rect 18880 29776 18932 29782
rect 18880 29718 18932 29724
rect 18892 29073 18920 29718
rect 18972 29708 19024 29714
rect 18972 29650 19024 29656
rect 18984 29306 19012 29650
rect 18972 29300 19024 29306
rect 18972 29242 19024 29248
rect 19076 29186 19104 30194
rect 19168 29646 19196 31282
rect 19524 31204 19576 31210
rect 19524 31146 19576 31152
rect 19340 31136 19392 31142
rect 19340 31078 19392 31084
rect 19246 30696 19302 30705
rect 19246 30631 19302 30640
rect 19156 29640 19208 29646
rect 19156 29582 19208 29588
rect 18984 29158 19104 29186
rect 19154 29200 19210 29209
rect 18878 29064 18934 29073
rect 18878 28999 18934 29008
rect 18984 28626 19012 29158
rect 19154 29135 19210 29144
rect 19168 28966 19196 29135
rect 19156 28960 19208 28966
rect 19156 28902 19208 28908
rect 19154 28792 19210 28801
rect 19076 28750 19154 28778
rect 18972 28620 19024 28626
rect 18972 28562 19024 28568
rect 18788 28212 18840 28218
rect 18788 28154 18840 28160
rect 18800 28082 18828 28154
rect 18788 28076 18840 28082
rect 18788 28018 18840 28024
rect 18708 27798 19012 27826
rect 18616 27662 18920 27690
rect 18524 27526 18736 27554
rect 18604 27464 18656 27470
rect 18604 27406 18656 27412
rect 18512 27396 18564 27402
rect 18512 27338 18564 27344
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18432 25974 18460 27270
rect 18524 27130 18552 27338
rect 18616 27130 18644 27406
rect 18512 27124 18564 27130
rect 18512 27066 18564 27072
rect 18604 27124 18656 27130
rect 18604 27066 18656 27072
rect 18512 26920 18564 26926
rect 18512 26862 18564 26868
rect 18420 25968 18472 25974
rect 18420 25910 18472 25916
rect 18328 25900 18380 25906
rect 18328 25842 18380 25848
rect 18420 25832 18472 25838
rect 18420 25774 18472 25780
rect 18144 25356 18196 25362
rect 18248 25350 18368 25378
rect 18144 25298 18196 25304
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 18248 24886 18276 25230
rect 18236 24880 18288 24886
rect 18236 24822 18288 24828
rect 17960 24676 18012 24682
rect 17960 24618 18012 24624
rect 17960 24336 18012 24342
rect 17682 24304 17738 24313
rect 17052 23718 17264 23746
rect 17328 24120 17356 24278
rect 17420 24262 17540 24290
rect 17512 24206 17540 24262
rect 17960 24278 18012 24284
rect 17682 24239 17738 24248
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17408 24132 17460 24138
rect 17328 24092 17408 24120
rect 16948 22160 17000 22166
rect 16948 22102 17000 22108
rect 17052 22030 17080 23718
rect 17328 23594 17356 24092
rect 17408 24074 17460 24080
rect 17696 23848 17724 24239
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17604 23820 17724 23848
rect 17500 23656 17552 23662
rect 17420 23616 17500 23644
rect 17316 23588 17368 23594
rect 17316 23530 17368 23536
rect 17328 23497 17356 23530
rect 17314 23488 17370 23497
rect 17314 23423 17370 23432
rect 17420 23118 17448 23616
rect 17500 23598 17552 23604
rect 17604 23526 17632 23820
rect 17776 23792 17828 23798
rect 17776 23734 17828 23740
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17696 23118 17724 23666
rect 17788 23526 17816 23734
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17684 23112 17736 23118
rect 17684 23054 17736 23060
rect 17144 22642 17172 23054
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17328 22642 17356 22986
rect 17132 22636 17184 22642
rect 17132 22578 17184 22584
rect 17316 22636 17368 22642
rect 17316 22578 17368 22584
rect 17224 22160 17276 22166
rect 17224 22102 17276 22108
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16960 21554 16988 21898
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 17052 21146 17080 21966
rect 17144 21690 17172 21966
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17236 21570 17264 22102
rect 17420 21690 17448 23054
rect 17500 22976 17552 22982
rect 17500 22918 17552 22924
rect 17512 22710 17540 22918
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 17500 22568 17552 22574
rect 17498 22536 17500 22545
rect 17552 22536 17554 22545
rect 17498 22471 17554 22480
rect 17592 21888 17644 21894
rect 17592 21830 17644 21836
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17132 21548 17184 21554
rect 17236 21542 17356 21570
rect 17132 21490 17184 21496
rect 17144 21434 17172 21490
rect 17144 21406 17264 21434
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 17144 21146 17172 21286
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17132 20936 17184 20942
rect 17236 20924 17264 21406
rect 17184 20896 17264 20924
rect 17132 20878 17184 20884
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16856 19848 16908 19854
rect 16960 19836 16988 20334
rect 16908 19808 16988 19836
rect 16856 19790 16908 19796
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16776 17678 16804 18702
rect 16856 18352 16908 18358
rect 16856 18294 16908 18300
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16776 17338 16804 17614
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16868 17116 16896 18294
rect 16960 18086 16988 19808
rect 17144 18698 17172 20878
rect 17222 20088 17278 20097
rect 17222 20023 17278 20032
rect 17236 19825 17264 20023
rect 17222 19816 17278 19825
rect 17222 19751 17278 19760
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17236 18970 17264 19110
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16960 17678 16988 18022
rect 17052 17728 17080 18226
rect 17224 17808 17276 17814
rect 17224 17750 17276 17756
rect 17052 17700 17172 17728
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16948 17128 17000 17134
rect 16868 17088 16948 17116
rect 16684 17054 16804 17082
rect 16948 17070 17000 17076
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16794 16712 16934
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16684 14414 16712 15846
rect 16776 15706 16804 17054
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16868 16250 16896 16526
rect 16960 16454 16988 17070
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16776 14414 16804 15506
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16684 13258 16712 14350
rect 16776 13954 16804 14350
rect 16868 14056 16896 15914
rect 16960 15570 16988 16390
rect 17052 16114 17080 17546
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 17144 15978 17172 17700
rect 17236 17270 17264 17750
rect 17328 17542 17356 21542
rect 17512 21078 17540 21626
rect 17500 21072 17552 21078
rect 17500 21014 17552 21020
rect 17408 20868 17460 20874
rect 17408 20810 17460 20816
rect 17420 19854 17448 20810
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17420 19378 17448 19790
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 17328 16658 17356 17478
rect 17512 16726 17540 21014
rect 17604 20806 17632 21830
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17604 18358 17632 20742
rect 17696 20058 17724 23054
rect 17788 23050 17816 23462
rect 17880 23118 17908 24142
rect 17972 23186 18000 24278
rect 18248 24206 18276 24822
rect 18340 24410 18368 25350
rect 18328 24404 18380 24410
rect 18328 24346 18380 24352
rect 18236 24200 18288 24206
rect 18236 24142 18288 24148
rect 17960 23180 18012 23186
rect 17960 23122 18012 23128
rect 17868 23112 17920 23118
rect 17868 23054 17920 23060
rect 17776 23044 17828 23050
rect 17776 22986 17828 22992
rect 17880 22642 17908 23054
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 17880 22166 17908 22578
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 17972 21026 18000 21490
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 17788 20998 18000 21026
rect 17788 20466 17816 20998
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17788 19990 17816 20198
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17880 19854 17908 20878
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17972 20058 18000 20402
rect 18064 20330 18092 21422
rect 18156 20641 18184 21422
rect 18248 21146 18276 24142
rect 18432 23594 18460 25774
rect 18524 25294 18552 26862
rect 18604 26580 18656 26586
rect 18604 26522 18656 26528
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 18524 24614 18552 25230
rect 18616 24954 18644 26522
rect 18708 25537 18736 27526
rect 18788 27328 18840 27334
rect 18788 27270 18840 27276
rect 18800 26353 18828 27270
rect 18892 26790 18920 27662
rect 18984 27606 19012 27798
rect 18972 27600 19024 27606
rect 18972 27542 19024 27548
rect 18984 27130 19012 27542
rect 18972 27124 19024 27130
rect 18972 27066 19024 27072
rect 18970 27024 19026 27033
rect 18970 26959 18972 26968
rect 19024 26959 19026 26968
rect 18972 26930 19024 26936
rect 18880 26784 18932 26790
rect 18880 26726 18932 26732
rect 18786 26344 18842 26353
rect 18786 26279 18842 26288
rect 18694 25528 18750 25537
rect 18694 25463 18750 25472
rect 18892 24954 18920 26726
rect 18970 26480 19026 26489
rect 18970 26415 19026 26424
rect 18984 25906 19012 26415
rect 18972 25900 19024 25906
rect 18972 25842 19024 25848
rect 19076 25702 19104 28750
rect 19154 28727 19210 28736
rect 19156 28144 19208 28150
rect 19156 28086 19208 28092
rect 19168 26586 19196 28086
rect 19156 26580 19208 26586
rect 19156 26522 19208 26528
rect 19260 26042 19288 30631
rect 19352 28490 19380 31078
rect 19536 30734 19564 31146
rect 19524 30728 19576 30734
rect 19524 30670 19576 30676
rect 19536 30598 19564 30670
rect 20088 30598 20116 35634
rect 20258 34368 20314 34377
rect 20258 34303 20314 34312
rect 20272 33998 20300 34303
rect 20260 33992 20312 33998
rect 20260 33934 20312 33940
rect 20272 33658 20300 33934
rect 20352 33856 20404 33862
rect 20352 33798 20404 33804
rect 20260 33652 20312 33658
rect 20260 33594 20312 33600
rect 20364 33522 20392 33798
rect 20352 33516 20404 33522
rect 20352 33458 20404 33464
rect 20168 33040 20220 33046
rect 20168 32982 20220 32988
rect 20180 31754 20208 32982
rect 20260 32904 20312 32910
rect 20260 32846 20312 32852
rect 20272 32502 20300 32846
rect 20260 32496 20312 32502
rect 20260 32438 20312 32444
rect 20352 31952 20404 31958
rect 20352 31894 20404 31900
rect 20180 31726 20300 31754
rect 20168 31680 20220 31686
rect 20168 31622 20220 31628
rect 19524 30592 19576 30598
rect 20076 30592 20128 30598
rect 19524 30534 19576 30540
rect 19996 30552 20076 30580
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19800 30388 19852 30394
rect 19800 30330 19852 30336
rect 19524 30320 19576 30326
rect 19524 30262 19576 30268
rect 19536 30025 19564 30262
rect 19522 30016 19578 30025
rect 19522 29951 19578 29960
rect 19706 29880 19762 29889
rect 19812 29850 19840 30330
rect 19996 30326 20024 30552
rect 20076 30534 20128 30540
rect 20074 30424 20130 30433
rect 20074 30359 20130 30368
rect 19984 30320 20036 30326
rect 19984 30262 20036 30268
rect 20088 30172 20116 30359
rect 19996 30144 20116 30172
rect 19892 30048 19944 30054
rect 19892 29990 19944 29996
rect 19706 29815 19762 29824
rect 19800 29844 19852 29850
rect 19720 29714 19748 29815
rect 19800 29786 19852 29792
rect 19904 29714 19932 29990
rect 19708 29708 19760 29714
rect 19708 29650 19760 29656
rect 19892 29708 19944 29714
rect 19892 29650 19944 29656
rect 19904 29492 19932 29650
rect 19444 29464 19932 29492
rect 19444 28994 19472 29464
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 19444 28966 19564 28994
rect 19904 28966 19932 29106
rect 19536 28529 19564 28966
rect 19892 28960 19944 28966
rect 19706 28928 19762 28937
rect 19628 28886 19706 28914
rect 19628 28626 19656 28886
rect 19892 28902 19944 28908
rect 19706 28863 19762 28872
rect 19904 28626 19932 28902
rect 19616 28620 19668 28626
rect 19616 28562 19668 28568
rect 19892 28620 19944 28626
rect 19892 28562 19944 28568
rect 19522 28520 19578 28529
rect 19340 28484 19392 28490
rect 19522 28455 19578 28464
rect 19340 28426 19392 28432
rect 19352 28014 19380 28426
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 19444 28200 19472 28358
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19444 28172 19564 28200
rect 19430 28112 19486 28121
rect 19430 28047 19486 28056
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19340 27464 19392 27470
rect 19340 27406 19392 27412
rect 19352 26926 19380 27406
rect 19444 27402 19472 28047
rect 19536 28014 19564 28172
rect 19628 28048 19932 28064
rect 19628 28042 19944 28048
rect 19628 28036 19892 28042
rect 19524 28008 19576 28014
rect 19524 27950 19576 27956
rect 19628 27946 19656 28036
rect 19892 27984 19944 27990
rect 19616 27940 19668 27946
rect 19616 27882 19668 27888
rect 19892 27872 19944 27878
rect 19892 27814 19944 27820
rect 19904 27402 19932 27814
rect 19432 27396 19484 27402
rect 19432 27338 19484 27344
rect 19892 27396 19944 27402
rect 19892 27338 19944 27344
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 19340 26920 19392 26926
rect 19340 26862 19392 26868
rect 19340 26784 19392 26790
rect 19340 26726 19392 26732
rect 19248 26036 19300 26042
rect 19248 25978 19300 25984
rect 19352 25906 19380 26726
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19064 25696 19116 25702
rect 19064 25638 19116 25644
rect 19156 25696 19208 25702
rect 19156 25638 19208 25644
rect 19340 25696 19392 25702
rect 19340 25638 19392 25644
rect 18604 24948 18656 24954
rect 18604 24890 18656 24896
rect 18880 24948 18932 24954
rect 18880 24890 18932 24896
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18420 23588 18472 23594
rect 18420 23530 18472 23536
rect 18524 22778 18552 24550
rect 18616 23746 18644 24890
rect 18696 24336 18748 24342
rect 18892 24324 18920 24890
rect 18748 24296 18920 24324
rect 18696 24278 18748 24284
rect 19076 24206 19104 25638
rect 19168 24410 19196 25638
rect 19248 25492 19300 25498
rect 19248 25434 19300 25440
rect 19156 24404 19208 24410
rect 19156 24346 19208 24352
rect 19154 24304 19210 24313
rect 19154 24239 19156 24248
rect 19208 24239 19210 24248
rect 19156 24210 19208 24216
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19260 24154 19288 25434
rect 19352 24682 19380 25638
rect 19340 24676 19392 24682
rect 19340 24618 19392 24624
rect 19444 24206 19472 26930
rect 19996 26790 20024 30144
rect 20180 30025 20208 31622
rect 20272 30977 20300 31726
rect 20258 30968 20314 30977
rect 20258 30903 20314 30912
rect 20364 30870 20392 31894
rect 20352 30864 20404 30870
rect 20352 30806 20404 30812
rect 20260 30728 20312 30734
rect 20260 30670 20312 30676
rect 20272 30161 20300 30670
rect 20364 30666 20392 30806
rect 20456 30734 20484 35702
rect 20548 34134 20576 36042
rect 20732 34950 20760 36654
rect 21008 35562 21036 37946
rect 22020 37874 22048 38150
rect 22468 38004 22520 38010
rect 22468 37946 22520 37952
rect 22744 38004 22796 38010
rect 22744 37946 22796 37952
rect 22008 37868 22060 37874
rect 22008 37810 22060 37816
rect 22020 37194 22048 37810
rect 22480 37738 22508 37946
rect 22652 37800 22704 37806
rect 22652 37742 22704 37748
rect 22468 37732 22520 37738
rect 22468 37674 22520 37680
rect 22376 37664 22428 37670
rect 22376 37606 22428 37612
rect 22388 37466 22416 37606
rect 22376 37460 22428 37466
rect 22376 37402 22428 37408
rect 22008 37188 22060 37194
rect 22008 37130 22060 37136
rect 22376 37120 22428 37126
rect 22376 37062 22428 37068
rect 22388 36922 22416 37062
rect 22376 36916 22428 36922
rect 22376 36858 22428 36864
rect 22468 36780 22520 36786
rect 22468 36722 22520 36728
rect 22480 36378 22508 36722
rect 22560 36644 22612 36650
rect 22560 36586 22612 36592
rect 22468 36372 22520 36378
rect 22468 36314 22520 36320
rect 22100 36236 22152 36242
rect 22100 36178 22152 36184
rect 21088 36100 21140 36106
rect 21088 36042 21140 36048
rect 20996 35556 21048 35562
rect 20996 35498 21048 35504
rect 21008 35154 21036 35498
rect 20996 35148 21048 35154
rect 20996 35090 21048 35096
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 20628 34400 20680 34406
rect 20628 34342 20680 34348
rect 20536 34128 20588 34134
rect 20536 34070 20588 34076
rect 20548 33998 20576 34070
rect 20640 33998 20668 34342
rect 20536 33992 20588 33998
rect 20536 33934 20588 33940
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20640 33640 20668 33934
rect 20548 33612 20668 33640
rect 20548 33318 20576 33612
rect 20628 33516 20680 33522
rect 20628 33458 20680 33464
rect 20640 33425 20668 33458
rect 20824 33454 20852 35022
rect 21008 34678 21036 35090
rect 20996 34672 21048 34678
rect 20996 34614 21048 34620
rect 21100 33658 21128 36042
rect 22112 35698 22140 36178
rect 22192 35760 22244 35766
rect 22192 35702 22244 35708
rect 21180 35692 21232 35698
rect 21180 35634 21232 35640
rect 22100 35692 22152 35698
rect 22100 35634 22152 35640
rect 21088 33652 21140 33658
rect 21088 33594 21140 33600
rect 21100 33561 21128 33594
rect 21086 33552 21142 33561
rect 21086 33487 21142 33496
rect 20812 33448 20864 33454
rect 20626 33416 20682 33425
rect 20864 33396 21036 33402
rect 20812 33390 21036 33396
rect 20824 33374 21036 33390
rect 20626 33351 20682 33360
rect 20536 33312 20588 33318
rect 20536 33254 20588 33260
rect 20626 33280 20682 33289
rect 20626 33215 20682 33224
rect 20536 33108 20588 33114
rect 20536 33050 20588 33056
rect 20548 32910 20576 33050
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20640 32008 20668 33215
rect 20904 32904 20956 32910
rect 20904 32846 20956 32852
rect 20720 32768 20772 32774
rect 20720 32710 20772 32716
rect 20548 31980 20668 32008
rect 20548 31754 20576 31980
rect 20628 31884 20680 31890
rect 20628 31826 20680 31832
rect 20536 31748 20588 31754
rect 20536 31690 20588 31696
rect 20548 31346 20576 31690
rect 20640 31346 20668 31826
rect 20732 31346 20760 32710
rect 20536 31340 20588 31346
rect 20536 31282 20588 31288
rect 20628 31340 20680 31346
rect 20628 31282 20680 31288
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20718 31104 20774 31113
rect 20916 31090 20944 32846
rect 20774 31062 20944 31090
rect 20718 31039 20774 31048
rect 20732 30870 20760 31039
rect 21008 30938 21036 33374
rect 21086 32872 21142 32881
rect 21086 32807 21142 32816
rect 21100 31346 21128 32807
rect 21192 31634 21220 35634
rect 21456 35624 21508 35630
rect 21456 35566 21508 35572
rect 21272 34672 21324 34678
rect 21272 34614 21324 34620
rect 21284 33658 21312 34614
rect 21272 33652 21324 33658
rect 21272 33594 21324 33600
rect 21468 33590 21496 35566
rect 22100 34672 22152 34678
rect 22020 34632 22100 34660
rect 21732 33992 21784 33998
rect 21730 33960 21732 33969
rect 21916 33992 21968 33998
rect 21784 33960 21786 33969
rect 21916 33934 21968 33940
rect 21730 33895 21786 33904
rect 21732 33856 21784 33862
rect 21732 33798 21784 33804
rect 21456 33584 21508 33590
rect 21508 33544 21588 33572
rect 21456 33526 21508 33532
rect 21456 33312 21508 33318
rect 21456 33254 21508 33260
rect 21468 32910 21496 33254
rect 21456 32904 21508 32910
rect 21456 32846 21508 32852
rect 21270 32464 21326 32473
rect 21270 32399 21272 32408
rect 21324 32399 21326 32408
rect 21364 32428 21416 32434
rect 21272 32370 21324 32376
rect 21364 32370 21416 32376
rect 21272 31816 21324 31822
rect 21270 31784 21272 31793
rect 21324 31784 21326 31793
rect 21270 31719 21326 31728
rect 21192 31606 21312 31634
rect 21180 31476 21232 31482
rect 21180 31418 21232 31424
rect 21088 31340 21140 31346
rect 21088 31282 21140 31288
rect 21192 31278 21220 31418
rect 21180 31272 21232 31278
rect 21180 31214 21232 31220
rect 20996 30932 21048 30938
rect 20996 30874 21048 30880
rect 20720 30864 20772 30870
rect 20720 30806 20772 30812
rect 20444 30728 20496 30734
rect 20444 30670 20496 30676
rect 20352 30660 20404 30666
rect 20352 30602 20404 30608
rect 20350 30560 20406 30569
rect 20350 30495 20406 30504
rect 20364 30394 20392 30495
rect 20352 30388 20404 30394
rect 20352 30330 20404 30336
rect 20258 30152 20314 30161
rect 20258 30087 20314 30096
rect 20352 30116 20404 30122
rect 20166 30016 20222 30025
rect 20166 29951 20222 29960
rect 20272 29866 20300 30087
rect 20352 30058 20404 30064
rect 20076 29844 20128 29850
rect 20076 29786 20128 29792
rect 20180 29838 20300 29866
rect 20088 28200 20116 29786
rect 20180 28422 20208 29838
rect 20258 29472 20314 29481
rect 20258 29407 20314 29416
rect 20272 28994 20300 29407
rect 20364 29238 20392 30058
rect 20456 30054 20484 30670
rect 20904 30592 20956 30598
rect 20904 30534 20956 30540
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20810 30288 20866 30297
rect 20534 30152 20590 30161
rect 20534 30087 20590 30096
rect 20548 30054 20576 30087
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 20536 30048 20588 30054
rect 20536 29990 20588 29996
rect 20640 29866 20668 30262
rect 20810 30223 20866 30232
rect 20824 30054 20852 30223
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20456 29838 20668 29866
rect 20720 29844 20772 29850
rect 20352 29232 20404 29238
rect 20352 29174 20404 29180
rect 20272 28966 20392 28994
rect 20260 28756 20312 28762
rect 20260 28698 20312 28704
rect 20272 28665 20300 28698
rect 20258 28656 20314 28665
rect 20258 28591 20314 28600
rect 20168 28416 20220 28422
rect 20168 28358 20220 28364
rect 20088 28172 20208 28200
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 19984 26784 20036 26790
rect 19984 26726 20036 26732
rect 20088 26353 20116 28018
rect 20180 27606 20208 28172
rect 20364 28098 20392 28966
rect 20272 28070 20392 28098
rect 20168 27600 20220 27606
rect 20168 27542 20220 27548
rect 20168 27328 20220 27334
rect 20168 27270 20220 27276
rect 20074 26344 20130 26353
rect 20180 26314 20208 27270
rect 20074 26279 20130 26288
rect 20168 26308 20220 26314
rect 20168 26250 20220 26256
rect 20076 26240 20128 26246
rect 20076 26182 20128 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19800 26036 19852 26042
rect 19800 25978 19852 25984
rect 19812 25906 19840 25978
rect 19892 25968 19944 25974
rect 19892 25910 19944 25916
rect 19800 25900 19852 25906
rect 19800 25842 19852 25848
rect 19524 25764 19576 25770
rect 19708 25764 19760 25770
rect 19576 25724 19708 25752
rect 19524 25706 19576 25712
rect 19708 25706 19760 25712
rect 19904 25158 19932 25910
rect 20088 25838 20116 26182
rect 20272 25974 20300 28070
rect 20352 28008 20404 28014
rect 20456 27996 20484 29838
rect 20720 29786 20772 29792
rect 20628 29776 20680 29782
rect 20628 29718 20680 29724
rect 20536 29640 20588 29646
rect 20536 29582 20588 29588
rect 20404 27968 20484 27996
rect 20352 27950 20404 27956
rect 20548 27962 20576 29582
rect 20640 29170 20668 29718
rect 20628 29164 20680 29170
rect 20628 29106 20680 29112
rect 20640 28558 20668 29106
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20732 28370 20760 29786
rect 20916 29492 20944 30534
rect 21088 30388 21140 30394
rect 21088 30330 21140 30336
rect 20996 29504 21048 29510
rect 20916 29464 20996 29492
rect 20996 29446 21048 29452
rect 20810 29336 20866 29345
rect 20994 29336 21050 29345
rect 20810 29271 20866 29280
rect 20916 29294 20994 29322
rect 20824 28558 20852 29271
rect 20916 29238 20944 29294
rect 20994 29271 21050 29280
rect 20904 29232 20956 29238
rect 20904 29174 20956 29180
rect 20812 28552 20864 28558
rect 20812 28494 20864 28500
rect 20732 28342 20852 28370
rect 20718 28248 20774 28257
rect 20718 28183 20774 28192
rect 20732 28150 20760 28183
rect 20720 28144 20772 28150
rect 20720 28086 20772 28092
rect 20260 25968 20312 25974
rect 20260 25910 20312 25916
rect 20076 25832 20128 25838
rect 20076 25774 20128 25780
rect 20258 25800 20314 25809
rect 20258 25735 20314 25744
rect 20272 25401 20300 25735
rect 20258 25392 20314 25401
rect 20258 25327 20314 25336
rect 20076 25220 20128 25226
rect 20076 25162 20128 25168
rect 19892 25152 19944 25158
rect 19892 25094 19944 25100
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 20088 24818 20116 25162
rect 19800 24812 19852 24818
rect 19800 24754 19852 24760
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19432 24200 19484 24206
rect 18708 23866 18736 24142
rect 19156 24132 19208 24138
rect 19260 24126 19380 24154
rect 19432 24142 19484 24148
rect 19156 24074 19208 24080
rect 19064 24064 19116 24070
rect 19064 24006 19116 24012
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18616 23718 18920 23746
rect 18602 23488 18658 23497
rect 18602 23423 18658 23432
rect 18616 23118 18644 23423
rect 18604 23112 18656 23118
rect 18604 23054 18656 23060
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 18800 21146 18828 22918
rect 18892 22094 18920 23718
rect 19076 22094 19104 24006
rect 19168 23730 19196 24074
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19260 23866 19288 24006
rect 19352 23866 19380 24126
rect 19536 24052 19564 24550
rect 19812 24274 19840 24754
rect 19800 24268 19852 24274
rect 19800 24210 19852 24216
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19444 24024 19564 24052
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19444 23746 19472 24024
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19708 23860 19760 23866
rect 19996 23848 20024 24142
rect 19708 23802 19760 23808
rect 19904 23820 20024 23848
rect 19352 23730 19472 23746
rect 19156 23724 19208 23730
rect 19156 23666 19208 23672
rect 19340 23724 19472 23730
rect 19392 23718 19472 23724
rect 19522 23760 19578 23769
rect 19522 23695 19524 23704
rect 19340 23666 19392 23672
rect 19576 23695 19578 23704
rect 19524 23666 19576 23672
rect 19352 22710 19380 23666
rect 19720 23050 19748 23802
rect 19904 23594 19932 23820
rect 19892 23588 19944 23594
rect 19892 23530 19944 23536
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 19812 23322 19840 23462
rect 19904 23322 19932 23530
rect 19800 23316 19852 23322
rect 19800 23258 19852 23264
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 19708 23044 19760 23050
rect 19708 22986 19760 22992
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 20088 22506 20116 24754
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 20180 23798 20208 24006
rect 20272 23798 20300 25327
rect 20364 25226 20392 27950
rect 20548 27934 20668 27962
rect 20536 27872 20588 27878
rect 20456 27820 20536 27826
rect 20456 27814 20588 27820
rect 20456 27798 20576 27814
rect 20456 27674 20484 27798
rect 20640 27690 20668 27934
rect 20444 27668 20496 27674
rect 20444 27610 20496 27616
rect 20548 27662 20668 27690
rect 20444 26308 20496 26314
rect 20444 26250 20496 26256
rect 20456 25906 20484 26250
rect 20548 25974 20576 27662
rect 20628 27600 20680 27606
rect 20628 27542 20680 27548
rect 20536 25968 20588 25974
rect 20536 25910 20588 25916
rect 20444 25900 20496 25906
rect 20444 25842 20496 25848
rect 20456 25498 20484 25842
rect 20444 25492 20496 25498
rect 20444 25434 20496 25440
rect 20640 25242 20668 27542
rect 20732 25294 20760 28086
rect 20824 26489 20852 28342
rect 20916 27985 20944 29174
rect 21100 29170 21128 30330
rect 21192 30326 21220 31214
rect 21284 30734 21312 31606
rect 21376 31482 21404 32370
rect 21468 31482 21496 32846
rect 21560 32774 21588 33544
rect 21548 32768 21600 32774
rect 21548 32710 21600 32716
rect 21364 31476 21416 31482
rect 21364 31418 21416 31424
rect 21456 31476 21508 31482
rect 21456 31418 21508 31424
rect 21468 31210 21496 31418
rect 21560 31249 21588 32710
rect 21640 32496 21692 32502
rect 21640 32438 21692 32444
rect 21652 31346 21680 32438
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 21744 31278 21772 33798
rect 21928 33658 21956 33934
rect 21916 33652 21968 33658
rect 21916 33594 21968 33600
rect 21822 33552 21878 33561
rect 21822 33487 21824 33496
rect 21876 33487 21878 33496
rect 21824 33458 21876 33464
rect 21836 31958 21864 33458
rect 21928 32910 21956 33594
rect 22020 33046 22048 34632
rect 22100 34614 22152 34620
rect 22100 34400 22152 34406
rect 22100 34342 22152 34348
rect 22112 33998 22140 34342
rect 22100 33992 22152 33998
rect 22100 33934 22152 33940
rect 22112 33318 22140 33934
rect 22100 33312 22152 33318
rect 22098 33280 22100 33289
rect 22152 33280 22154 33289
rect 22098 33215 22154 33224
rect 22008 33040 22060 33046
rect 22204 32994 22232 35702
rect 22572 35698 22600 36586
rect 22284 35692 22336 35698
rect 22284 35634 22336 35640
rect 22376 35692 22428 35698
rect 22376 35634 22428 35640
rect 22560 35692 22612 35698
rect 22560 35634 22612 35640
rect 22296 34950 22324 35634
rect 22284 34944 22336 34950
rect 22284 34886 22336 34892
rect 22296 34610 22324 34886
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 22284 34400 22336 34406
rect 22284 34342 22336 34348
rect 22296 33998 22324 34342
rect 22284 33992 22336 33998
rect 22284 33934 22336 33940
rect 22008 32982 22060 32988
rect 22112 32966 22232 32994
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 22008 32020 22060 32026
rect 22008 31962 22060 31968
rect 21824 31952 21876 31958
rect 21824 31894 21876 31900
rect 22020 31822 22048 31962
rect 22112 31822 22140 32966
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 22204 32230 22232 32846
rect 22284 32428 22336 32434
rect 22284 32370 22336 32376
rect 22192 32224 22244 32230
rect 22192 32166 22244 32172
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 21822 31512 21878 31521
rect 21822 31447 21878 31456
rect 21836 31346 21864 31447
rect 21824 31340 21876 31346
rect 21824 31282 21876 31288
rect 21732 31272 21784 31278
rect 21546 31240 21602 31249
rect 21456 31204 21508 31210
rect 21732 31214 21784 31220
rect 21546 31175 21548 31184
rect 21456 31146 21508 31152
rect 21600 31175 21602 31184
rect 21548 31146 21600 31152
rect 21468 31090 21496 31146
rect 21468 31062 21588 31090
rect 21362 30968 21418 30977
rect 21362 30903 21418 30912
rect 21376 30734 21404 30903
rect 21272 30728 21324 30734
rect 21272 30670 21324 30676
rect 21364 30728 21416 30734
rect 21364 30670 21416 30676
rect 21180 30320 21232 30326
rect 21180 30262 21232 30268
rect 21284 29850 21312 30670
rect 21272 29844 21324 29850
rect 21272 29786 21324 29792
rect 21284 29646 21312 29786
rect 21272 29640 21324 29646
rect 21272 29582 21324 29588
rect 21088 29164 21140 29170
rect 21376 29152 21404 30670
rect 21560 30122 21588 31062
rect 21548 30116 21600 30122
rect 21548 30058 21600 30064
rect 21640 29708 21692 29714
rect 21640 29650 21692 29656
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 21468 29306 21496 29582
rect 21546 29472 21602 29481
rect 21546 29407 21602 29416
rect 21456 29300 21508 29306
rect 21456 29242 21508 29248
rect 21376 29124 21496 29152
rect 21088 29106 21140 29112
rect 21468 29050 21496 29124
rect 21376 29022 21496 29050
rect 21272 29006 21324 29012
rect 21272 28948 21324 28954
rect 21284 28558 21312 28948
rect 20996 28552 21048 28558
rect 20996 28494 21048 28500
rect 21272 28552 21324 28558
rect 21272 28494 21324 28500
rect 20902 27976 20958 27985
rect 20902 27911 20958 27920
rect 20810 26480 20866 26489
rect 20810 26415 20866 26424
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 20824 26042 20852 26318
rect 20812 26036 20864 26042
rect 20812 25978 20864 25984
rect 20916 25702 20944 26318
rect 21008 25906 21036 28494
rect 21088 28416 21140 28422
rect 21088 28358 21140 28364
rect 21100 27402 21128 28358
rect 21272 27872 21324 27878
rect 21178 27840 21234 27849
rect 21272 27814 21324 27820
rect 21178 27775 21234 27784
rect 21088 27396 21140 27402
rect 21088 27338 21140 27344
rect 21192 26042 21220 27775
rect 21284 27538 21312 27814
rect 21272 27532 21324 27538
rect 21272 27474 21324 27480
rect 21180 26036 21232 26042
rect 21180 25978 21232 25984
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 20904 25696 20956 25702
rect 20904 25638 20956 25644
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 20916 25430 20944 25638
rect 20904 25424 20956 25430
rect 20904 25366 20956 25372
rect 21008 25362 21036 25638
rect 20996 25356 21048 25362
rect 20996 25298 21048 25304
rect 20352 25220 20404 25226
rect 20352 25162 20404 25168
rect 20548 25214 20668 25242
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20444 24744 20496 24750
rect 20444 24686 20496 24692
rect 20352 24336 20404 24342
rect 20352 24278 20404 24284
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 20260 23792 20312 23798
rect 20260 23734 20312 23740
rect 20364 23594 20392 24278
rect 20456 24206 20484 24686
rect 20548 24206 20576 25214
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20536 24200 20588 24206
rect 20536 24142 20588 24148
rect 20456 23610 20484 24142
rect 20548 23866 20576 24142
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 20352 23588 20404 23594
rect 20456 23582 20576 23610
rect 20352 23530 20404 23536
rect 20364 23100 20392 23530
rect 20548 23186 20576 23582
rect 20536 23180 20588 23186
rect 20536 23122 20588 23128
rect 20640 23118 20668 25094
rect 21100 24886 21128 25638
rect 21192 25294 21220 25978
rect 21272 25696 21324 25702
rect 21272 25638 21324 25644
rect 21284 25430 21312 25638
rect 21272 25424 21324 25430
rect 21272 25366 21324 25372
rect 21180 25288 21232 25294
rect 21180 25230 21232 25236
rect 21180 25152 21232 25158
rect 21180 25094 21232 25100
rect 20996 24880 21048 24886
rect 20996 24822 21048 24828
rect 21088 24880 21140 24886
rect 21088 24822 21140 24828
rect 21008 24732 21036 24822
rect 21192 24732 21220 25094
rect 21008 24704 21220 24732
rect 21284 24614 21312 25366
rect 21376 24614 21404 29022
rect 21454 28928 21510 28937
rect 21454 28863 21510 28872
rect 21468 28082 21496 28863
rect 21560 28422 21588 29407
rect 21652 29306 21680 29650
rect 21640 29300 21692 29306
rect 21640 29242 21692 29248
rect 21638 29200 21694 29209
rect 21638 29135 21640 29144
rect 21692 29135 21694 29144
rect 21640 29106 21692 29112
rect 21640 28552 21692 28558
rect 21640 28494 21692 28500
rect 21548 28416 21600 28422
rect 21548 28358 21600 28364
rect 21456 28076 21508 28082
rect 21456 28018 21508 28024
rect 21456 27396 21508 27402
rect 21456 27338 21508 27344
rect 21468 26194 21496 27338
rect 21560 26314 21588 28358
rect 21652 28082 21680 28494
rect 21640 28076 21692 28082
rect 21640 28018 21692 28024
rect 21744 27538 21772 31214
rect 21928 30938 21956 31758
rect 21916 30932 21968 30938
rect 21916 30874 21968 30880
rect 22008 30252 22060 30258
rect 22008 30194 22060 30200
rect 22020 29850 22048 30194
rect 22008 29844 22060 29850
rect 22008 29786 22060 29792
rect 21824 29504 21876 29510
rect 21824 29446 21876 29452
rect 21836 29170 21864 29446
rect 22112 29170 22140 31758
rect 22204 31482 22232 32166
rect 22192 31476 22244 31482
rect 22192 31418 22244 31424
rect 22296 31362 22324 32370
rect 22388 31822 22416 35634
rect 22560 35148 22612 35154
rect 22560 35090 22612 35096
rect 22572 34746 22600 35090
rect 22560 34740 22612 34746
rect 22560 34682 22612 34688
rect 22558 34232 22614 34241
rect 22558 34167 22614 34176
rect 22468 33992 22520 33998
rect 22468 33934 22520 33940
rect 22480 33862 22508 33934
rect 22572 33862 22600 34167
rect 22468 33856 22520 33862
rect 22466 33824 22468 33833
rect 22560 33856 22612 33862
rect 22520 33824 22522 33833
rect 22560 33798 22612 33804
rect 22466 33759 22522 33768
rect 22664 33658 22692 37742
rect 22756 37262 22784 37946
rect 23112 37868 23164 37874
rect 23112 37810 23164 37816
rect 23664 37868 23716 37874
rect 23664 37810 23716 37816
rect 23756 37868 23808 37874
rect 23756 37810 23808 37816
rect 22926 37360 22982 37369
rect 22926 37295 22928 37304
rect 22980 37295 22982 37304
rect 22928 37266 22980 37272
rect 22744 37256 22796 37262
rect 22744 37198 22796 37204
rect 22836 37188 22888 37194
rect 22836 37130 22888 37136
rect 22848 36174 22876 37130
rect 23020 36372 23072 36378
rect 23020 36314 23072 36320
rect 22836 36168 22888 36174
rect 22836 36110 22888 36116
rect 22928 36032 22980 36038
rect 22928 35974 22980 35980
rect 22940 35698 22968 35974
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22928 35692 22980 35698
rect 22928 35634 22980 35640
rect 22744 35624 22796 35630
rect 22744 35566 22796 35572
rect 22468 33652 22520 33658
rect 22468 33594 22520 33600
rect 22652 33652 22704 33658
rect 22652 33594 22704 33600
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22204 31334 22324 31362
rect 22204 29458 22232 31334
rect 22284 30116 22336 30122
rect 22284 30058 22336 30064
rect 22296 29578 22324 30058
rect 22284 29572 22336 29578
rect 22284 29514 22336 29520
rect 22204 29430 22324 29458
rect 21824 29164 21876 29170
rect 21824 29106 21876 29112
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 22192 29164 22244 29170
rect 22192 29106 22244 29112
rect 22020 28558 22048 29106
rect 22112 29073 22140 29106
rect 22098 29064 22154 29073
rect 22098 28999 22154 29008
rect 22008 28552 22060 28558
rect 22008 28494 22060 28500
rect 22204 28150 22232 29106
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 21824 28008 21876 28014
rect 21824 27950 21876 27956
rect 21916 28008 21968 28014
rect 21916 27950 21968 27956
rect 21732 27532 21784 27538
rect 21732 27474 21784 27480
rect 21548 26308 21600 26314
rect 21548 26250 21600 26256
rect 21468 26166 21588 26194
rect 21454 25800 21510 25809
rect 21454 25735 21510 25744
rect 21468 25294 21496 25735
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21560 24818 21588 26166
rect 21744 25294 21772 27474
rect 21836 26489 21864 27950
rect 21928 27713 21956 27950
rect 21914 27704 21970 27713
rect 21914 27639 21970 27648
rect 22204 27334 22232 28086
rect 22296 27878 22324 29430
rect 22388 29238 22416 31758
rect 22376 29232 22428 29238
rect 22376 29174 22428 29180
rect 22376 28552 22428 28558
rect 22376 28494 22428 28500
rect 22284 27872 22336 27878
rect 22284 27814 22336 27820
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 22192 27124 22244 27130
rect 22192 27066 22244 27072
rect 21822 26480 21878 26489
rect 21822 26415 21878 26424
rect 22204 25906 22232 27066
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22296 25786 22324 27814
rect 22388 25922 22416 28494
rect 22480 26042 22508 33594
rect 22560 32020 22612 32026
rect 22560 31962 22612 31968
rect 22572 31929 22600 31962
rect 22756 31958 22784 35566
rect 22848 33658 22876 35634
rect 22928 34944 22980 34950
rect 22928 34886 22980 34892
rect 22940 33969 22968 34886
rect 23032 34746 23060 36314
rect 23020 34740 23072 34746
rect 23020 34682 23072 34688
rect 23124 34610 23152 37810
rect 23480 37324 23532 37330
rect 23480 37266 23532 37272
rect 23296 37256 23348 37262
rect 23296 37198 23348 37204
rect 23308 36242 23336 37198
rect 23492 36786 23520 37266
rect 23572 37188 23624 37194
rect 23572 37130 23624 37136
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23480 36644 23532 36650
rect 23480 36586 23532 36592
rect 23492 36258 23520 36586
rect 23584 36378 23612 37130
rect 23572 36372 23624 36378
rect 23572 36314 23624 36320
rect 23296 36236 23348 36242
rect 23492 36230 23612 36258
rect 23296 36178 23348 36184
rect 23204 36168 23256 36174
rect 23204 36110 23256 36116
rect 23216 35766 23244 36110
rect 23296 35828 23348 35834
rect 23296 35770 23348 35776
rect 23204 35760 23256 35766
rect 23204 35702 23256 35708
rect 23216 34678 23244 35702
rect 23204 34672 23256 34678
rect 23204 34614 23256 34620
rect 23112 34604 23164 34610
rect 23112 34546 23164 34552
rect 23020 34400 23072 34406
rect 23020 34342 23072 34348
rect 23032 34105 23060 34342
rect 23018 34096 23074 34105
rect 23018 34031 23074 34040
rect 22926 33960 22982 33969
rect 22926 33895 22982 33904
rect 22836 33652 22888 33658
rect 22836 33594 22888 33600
rect 22836 32904 22888 32910
rect 22834 32872 22836 32881
rect 22888 32872 22890 32881
rect 22834 32807 22890 32816
rect 22848 32502 22876 32807
rect 22836 32496 22888 32502
rect 22836 32438 22888 32444
rect 22836 32224 22888 32230
rect 22836 32166 22888 32172
rect 22744 31952 22796 31958
rect 22558 31920 22614 31929
rect 22744 31894 22796 31900
rect 22558 31855 22614 31864
rect 22560 31680 22612 31686
rect 22560 31622 22612 31628
rect 22652 31680 22704 31686
rect 22652 31622 22704 31628
rect 22744 31680 22796 31686
rect 22744 31622 22796 31628
rect 22572 31346 22600 31622
rect 22560 31340 22612 31346
rect 22560 31282 22612 31288
rect 22560 30864 22612 30870
rect 22560 30806 22612 30812
rect 22572 29170 22600 30806
rect 22664 30326 22692 31622
rect 22756 31385 22784 31622
rect 22742 31376 22798 31385
rect 22848 31346 22876 32166
rect 22940 31754 22968 33895
rect 23032 33862 23060 34031
rect 23204 33992 23256 33998
rect 23110 33960 23166 33969
rect 23204 33934 23256 33940
rect 23110 33895 23166 33904
rect 23124 33862 23152 33895
rect 23020 33856 23072 33862
rect 23020 33798 23072 33804
rect 23112 33856 23164 33862
rect 23216 33833 23244 33934
rect 23112 33798 23164 33804
rect 23202 33824 23258 33833
rect 23202 33759 23258 33768
rect 23032 33658 23244 33674
rect 23020 33652 23244 33658
rect 23072 33646 23244 33652
rect 23020 33594 23072 33600
rect 23112 32360 23164 32366
rect 23112 32302 23164 32308
rect 23124 31958 23152 32302
rect 23020 31952 23072 31958
rect 23020 31894 23072 31900
rect 23112 31952 23164 31958
rect 23112 31894 23164 31900
rect 23032 31804 23060 31894
rect 23112 31816 23164 31822
rect 23032 31776 23112 31804
rect 23112 31758 23164 31764
rect 22928 31748 22980 31754
rect 22928 31690 22980 31696
rect 22742 31311 22798 31320
rect 22836 31340 22888 31346
rect 22836 31282 22888 31288
rect 22940 30546 22968 31690
rect 23018 31376 23074 31385
rect 23018 31311 23020 31320
rect 23072 31311 23074 31320
rect 23020 31282 23072 31288
rect 23020 31136 23072 31142
rect 23020 31078 23072 31084
rect 22756 30518 22968 30546
rect 22652 30320 22704 30326
rect 22652 30262 22704 30268
rect 22756 29646 22784 30518
rect 22834 30424 22890 30433
rect 22834 30359 22890 30368
rect 22744 29640 22796 29646
rect 22742 29608 22744 29617
rect 22796 29608 22798 29617
rect 22742 29543 22798 29552
rect 22652 29504 22704 29510
rect 22652 29446 22704 29452
rect 22664 29170 22692 29446
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22558 28656 22614 28665
rect 22558 28591 22614 28600
rect 22572 28558 22600 28591
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22572 26790 22600 28494
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 22652 26512 22704 26518
rect 22652 26454 22704 26460
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22388 25894 22508 25922
rect 22664 25906 22692 26454
rect 22756 26246 22784 26930
rect 22744 26240 22796 26246
rect 22744 26182 22796 26188
rect 21928 25758 22324 25786
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 21744 24818 21772 25230
rect 21548 24812 21600 24818
rect 21548 24754 21600 24760
rect 21732 24812 21784 24818
rect 21732 24754 21784 24760
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21364 24608 21416 24614
rect 21364 24550 21416 24556
rect 21376 23798 21404 24550
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21730 23760 21786 23769
rect 20812 23724 20864 23730
rect 21928 23746 21956 25758
rect 22284 25696 22336 25702
rect 22284 25638 22336 25644
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22192 25288 22244 25294
rect 22192 25230 22244 25236
rect 22008 25220 22060 25226
rect 22008 25162 22060 25168
rect 22020 24886 22048 25162
rect 22008 24880 22060 24886
rect 22008 24822 22060 24828
rect 22020 24274 22048 24822
rect 22204 24750 22232 25230
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 22100 24336 22152 24342
rect 22100 24278 22152 24284
rect 22008 24268 22060 24274
rect 22008 24210 22060 24216
rect 22112 24177 22140 24278
rect 22098 24168 22154 24177
rect 22098 24103 22154 24112
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 21786 23718 21956 23746
rect 21730 23695 21786 23704
rect 20812 23666 20864 23672
rect 20824 23322 20852 23666
rect 22204 23594 22232 24006
rect 22192 23588 22244 23594
rect 22192 23530 22244 23536
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 22192 23180 22244 23186
rect 22192 23122 22244 23128
rect 20444 23112 20496 23118
rect 20364 23072 20444 23100
rect 20444 23054 20496 23060
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20260 23044 20312 23050
rect 20260 22986 20312 22992
rect 19248 22500 19300 22506
rect 19248 22442 19300 22448
rect 20076 22500 20128 22506
rect 20076 22442 20128 22448
rect 19260 22166 19288 22442
rect 19248 22160 19300 22166
rect 19248 22102 19300 22108
rect 18892 22066 19012 22094
rect 19076 22066 19196 22094
rect 18984 21690 19012 22066
rect 18972 21684 19024 21690
rect 18972 21626 19024 21632
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18236 21140 18288 21146
rect 18512 21140 18564 21146
rect 18236 21082 18288 21088
rect 18340 21100 18512 21128
rect 18142 20632 18198 20641
rect 18142 20567 18198 20576
rect 18156 20466 18184 20567
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18052 20324 18104 20330
rect 18052 20266 18104 20272
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17880 19360 17908 19790
rect 17972 19718 18000 19994
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17880 19332 18000 19360
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17592 18352 17644 18358
rect 17592 18294 17644 18300
rect 17696 17678 17724 18702
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17788 17610 17816 19246
rect 17972 18086 18000 19332
rect 18064 18970 18092 20266
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18248 19786 18276 19994
rect 18236 19780 18288 19786
rect 18236 19722 18288 19728
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18156 19514 18184 19654
rect 18144 19508 18196 19514
rect 18144 19450 18196 19456
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18052 18760 18104 18766
rect 18050 18728 18052 18737
rect 18104 18728 18106 18737
rect 18050 18663 18106 18672
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 18064 17678 18092 18566
rect 18156 17678 18184 19450
rect 18248 18290 18276 19722
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18248 18193 18276 18226
rect 18234 18184 18290 18193
rect 18234 18119 18290 18128
rect 18234 17912 18290 17921
rect 18234 17847 18290 17856
rect 18248 17678 18276 17847
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 18340 17202 18368 21100
rect 18512 21082 18564 21088
rect 18788 21140 18840 21146
rect 18788 21082 18840 21088
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18524 20466 18552 20742
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18616 20466 18644 20538
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18604 20460 18656 20466
rect 18800 20448 18828 20878
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18656 20420 18828 20448
rect 18604 20402 18656 20408
rect 18432 18766 18460 20402
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18616 18902 18644 20198
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 18708 19854 18736 19994
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18604 18896 18656 18902
rect 18604 18838 18656 18844
rect 18420 18760 18472 18766
rect 18418 18728 18420 18737
rect 18472 18728 18474 18737
rect 18418 18663 18474 18672
rect 18432 18358 18460 18663
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18418 17912 18474 17921
rect 18418 17847 18474 17856
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 17500 16720 17552 16726
rect 17420 16680 17500 16708
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17328 16250 17356 16594
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 17132 15972 17184 15978
rect 17132 15914 17184 15920
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 16960 14346 16988 14962
rect 17052 14618 17080 14962
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 16948 14068 17000 14074
rect 16868 14028 16948 14056
rect 16948 14010 17000 14016
rect 16776 13926 16896 13954
rect 17144 13938 17172 15914
rect 17236 15026 17264 16118
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 16868 13870 16896 13926
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 15948 9438 16068 9466
rect 16316 12838 16528 12866
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15672 7954 15700 8230
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15580 7002 15608 7142
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15764 6866 15792 8910
rect 15948 8906 15976 9438
rect 16316 9382 16344 12838
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16408 12374 16436 12582
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16500 11014 16528 12174
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16500 10674 16528 10950
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16500 9704 16528 10610
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16500 9676 16620 9704
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16040 8906 16068 9318
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 16028 8900 16080 8906
rect 16592 8888 16620 9676
rect 16684 9586 16712 9862
rect 16776 9674 16804 13466
rect 16868 13462 16896 13806
rect 17236 13530 17264 14962
rect 17328 14006 17356 16186
rect 17420 14618 17448 16680
rect 17500 16662 17552 16668
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17604 15609 17632 16526
rect 17684 15632 17736 15638
rect 17590 15600 17646 15609
rect 17684 15574 17736 15580
rect 17590 15535 17646 15544
rect 17696 15026 17724 15574
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17696 14482 17724 14758
rect 17776 14544 17828 14550
rect 17774 14512 17776 14521
rect 17828 14512 17830 14521
rect 17684 14476 17736 14482
rect 17774 14447 17830 14456
rect 17684 14418 17736 14424
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 17420 13938 17448 14282
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17880 13734 17908 17138
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 17972 15570 18000 16526
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18156 16114 18184 16390
rect 18248 16114 18276 16934
rect 18432 16658 18460 17847
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18524 16454 18552 18022
rect 18616 17678 18644 18838
rect 18800 18714 18828 20420
rect 18892 19718 18920 20538
rect 18984 19836 19012 21422
rect 19062 20632 19118 20641
rect 19062 20567 19118 20576
rect 19076 20398 19104 20567
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19064 19848 19116 19854
rect 18984 19808 19064 19836
rect 19064 19790 19116 19796
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 18696 18692 18748 18698
rect 18800 18686 18920 18714
rect 18696 18634 18748 18640
rect 18708 17678 18736 18634
rect 18892 18630 18920 18686
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 18800 17678 18828 18566
rect 18892 18086 18920 18566
rect 18984 18290 19012 18906
rect 19064 18352 19116 18358
rect 19062 18320 19064 18329
rect 19116 18320 19118 18329
rect 18972 18284 19024 18290
rect 19062 18255 19118 18264
rect 18972 18226 19024 18232
rect 18970 18184 19026 18193
rect 19026 18142 19104 18170
rect 18970 18119 19026 18128
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 16590 18644 17478
rect 18708 16998 18736 17614
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18892 16114 18920 17478
rect 18984 17202 19012 17478
rect 19076 17338 19104 18142
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 19064 16516 19116 16522
rect 19064 16458 19116 16464
rect 19076 16250 19104 16458
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18340 15910 18368 16050
rect 18328 15904 18380 15910
rect 18328 15846 18380 15852
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18616 15570 18644 15846
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 18248 14958 18276 15370
rect 18616 15026 18644 15506
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16868 12442 16896 12786
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16776 9646 16896 9674
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16764 8900 16816 8906
rect 16592 8860 16764 8888
rect 16028 8842 16080 8848
rect 16764 8842 16816 8848
rect 16776 8498 16804 8842
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15396 6202 15424 6258
rect 15396 6174 15516 6202
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15212 5710 15240 6054
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15212 5370 15240 5646
rect 15396 5574 15424 6054
rect 15488 5914 15516 6174
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15764 5778 15792 6802
rect 16776 6730 16804 8434
rect 16868 7818 16896 9646
rect 16960 9518 16988 10610
rect 17052 10470 17080 10950
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 17144 10266 17172 10610
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 17328 8566 17356 9522
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17420 8498 17448 13670
rect 17880 13530 17908 13670
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17592 11620 17644 11626
rect 17696 11608 17724 12038
rect 17644 11580 17724 11608
rect 17592 11562 17644 11568
rect 17604 11354 17632 11562
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17498 10568 17554 10577
rect 17498 10503 17500 10512
rect 17552 10503 17554 10512
rect 17500 10474 17552 10480
rect 17788 9674 17816 12242
rect 18248 12238 18276 14894
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18432 13530 18460 13738
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18708 13326 18736 15846
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18972 15632 19024 15638
rect 18972 15574 19024 15580
rect 18788 15428 18840 15434
rect 18788 15370 18840 15376
rect 18800 15162 18828 15370
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18696 13320 18748 13326
rect 18524 13280 18696 13308
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 18340 12442 18368 13194
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18328 12300 18380 12306
rect 18524 12288 18552 13280
rect 18696 13262 18748 13268
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18708 13025 18736 13126
rect 18694 13016 18750 13025
rect 18694 12951 18750 12960
rect 18380 12260 18552 12288
rect 18328 12242 18380 12248
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18248 11150 18276 12174
rect 18694 11656 18750 11665
rect 18694 11591 18696 11600
rect 18748 11591 18750 11600
rect 18696 11562 18748 11568
rect 18800 11286 18828 14826
rect 18892 11830 18920 15574
rect 18984 15366 19012 15574
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18984 12238 19012 15302
rect 19168 13802 19196 22066
rect 19248 22024 19300 22030
rect 19984 22024 20036 22030
rect 19248 21966 19300 21972
rect 19260 21554 19288 21966
rect 19352 21962 19932 21978
rect 19984 21966 20036 21972
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 19340 21956 19944 21962
rect 19392 21950 19892 21956
rect 19340 21898 19392 21904
rect 19892 21898 19944 21904
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19340 21616 19392 21622
rect 19340 21558 19392 21564
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19352 21434 19380 21558
rect 19444 21486 19472 21830
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21486 20024 21966
rect 20074 21856 20130 21865
rect 20074 21791 20130 21800
rect 20088 21690 20116 21791
rect 20180 21690 20208 21966
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 19260 21406 19380 21434
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19260 20466 19288 21406
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19352 20262 19380 20742
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19260 19446 19288 19722
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 19260 18766 19288 19382
rect 19352 19378 19380 20198
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19444 18970 19472 21422
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19892 20256 19944 20262
rect 19996 20244 20024 20878
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 19944 20216 20024 20244
rect 19892 20198 19944 20204
rect 19904 19854 19932 20198
rect 20088 19922 20116 20402
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19984 19848 20036 19854
rect 20180 19802 20208 20198
rect 19984 19790 20036 19796
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 19514 20024 19790
rect 20088 19774 20208 19802
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19260 18086 19288 18702
rect 19352 18426 19380 18770
rect 19536 18766 19564 19450
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19628 18766 19656 19314
rect 19996 18970 20024 19314
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19996 18834 20024 18906
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19616 18760 19668 18766
rect 19668 18720 19840 18748
rect 19616 18702 19668 18708
rect 19812 18714 19840 18720
rect 19812 18686 20024 18714
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19352 17678 19380 18362
rect 19996 18358 20024 18686
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 19616 18284 19668 18290
rect 19616 18226 19668 18232
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19444 17678 19472 18158
rect 19628 18086 19656 18226
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19352 16561 19380 16730
rect 19338 16552 19394 16561
rect 19338 16487 19394 16496
rect 19352 15366 19380 16487
rect 19444 16250 19472 17274
rect 19720 17202 19748 17274
rect 19996 17270 20024 17614
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19628 16980 19656 17138
rect 19800 16992 19852 16998
rect 19628 16952 19800 16980
rect 19800 16934 19852 16940
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19444 15026 19472 15438
rect 20088 15434 20116 19774
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20180 19310 20208 19654
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 20180 18970 20208 19246
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 20180 17270 20208 17614
rect 20168 17264 20220 17270
rect 20168 17206 20220 17212
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19996 15026 20024 15302
rect 20180 15026 20208 17070
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19156 13796 19208 13802
rect 19156 13738 19208 13744
rect 19168 13258 19196 13738
rect 19352 13546 19380 14214
rect 19444 14074 19472 14826
rect 19996 14278 20024 14962
rect 20180 14550 20208 14962
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19260 13518 19380 13546
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19260 12918 19288 13518
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 18788 11280 18840 11286
rect 18788 11222 18840 11228
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18248 10674 18276 11086
rect 18800 10674 18828 11222
rect 18892 10810 18920 11766
rect 19260 11558 19288 12378
rect 19352 12238 19380 13398
rect 19444 12646 19472 13670
rect 19628 13326 19656 13874
rect 19720 13530 19748 13874
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19996 12782 20024 14214
rect 20088 14006 20116 14350
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20088 12986 20116 13262
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20180 12850 20208 13126
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19904 12374 19932 12582
rect 19892 12368 19944 12374
rect 19892 12310 19944 12316
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19260 11286 19288 11494
rect 19444 11354 19472 12038
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18234 10432 18290 10441
rect 18064 10062 18092 10406
rect 18234 10367 18290 10376
rect 18248 10062 18276 10367
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 17604 9646 17816 9674
rect 18064 9654 18092 9998
rect 18052 9648 18104 9654
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17512 8498 17540 9454
rect 17604 9042 17632 9646
rect 18052 9590 18104 9596
rect 18340 9586 18368 9998
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18248 9178 18276 9454
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18340 9178 18368 9386
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15396 5166 15424 5510
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15856 4826 15884 5102
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15948 4622 15976 5578
rect 16132 5234 16160 5578
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 16316 4622 16344 5850
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16408 4826 16436 4966
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16500 4622 16528 6054
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16684 4826 16712 5102
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16776 4486 16804 6666
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17144 5370 17172 5646
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 17236 3194 17264 8298
rect 17604 7886 17632 8978
rect 18432 8634 18460 9998
rect 18708 8974 18736 10202
rect 18800 10062 18828 10610
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18892 8498 18920 10746
rect 19260 10266 19288 11222
rect 20088 11150 20116 12106
rect 20272 11286 20300 22986
rect 20456 22778 20484 23054
rect 20444 22772 20496 22778
rect 22204 22760 22232 23122
rect 22296 23118 22324 25638
rect 22388 25294 22416 25638
rect 22480 25498 22508 25894
rect 22652 25900 22704 25906
rect 22652 25842 22704 25848
rect 22560 25764 22612 25770
rect 22560 25706 22612 25712
rect 22572 25498 22600 25706
rect 22468 25492 22520 25498
rect 22468 25434 22520 25440
rect 22560 25492 22612 25498
rect 22560 25434 22612 25440
rect 22652 25424 22704 25430
rect 22652 25366 22704 25372
rect 22376 25288 22428 25294
rect 22664 25242 22692 25366
rect 22376 25230 22428 25236
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22204 22732 22324 22760
rect 20444 22714 20496 22720
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20364 21690 20392 21898
rect 20352 21684 20404 21690
rect 20404 21644 20484 21672
rect 20352 21626 20404 21632
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20364 21146 20392 21490
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20364 20942 20392 21082
rect 20456 20942 20484 21644
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20444 20936 20496 20942
rect 20496 20896 20668 20924
rect 20444 20878 20496 20884
rect 20352 20800 20404 20806
rect 20350 20768 20352 20777
rect 20444 20800 20496 20806
rect 20404 20768 20406 20777
rect 20444 20742 20496 20748
rect 20350 20703 20406 20712
rect 20364 20466 20392 20703
rect 20456 20602 20484 20742
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20364 19854 20392 20198
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20456 18290 20484 20538
rect 20640 20466 20668 20896
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20548 19378 20576 19790
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20640 18766 20668 19654
rect 20732 18970 20760 22578
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21180 21616 21232 21622
rect 21180 21558 21232 21564
rect 20994 21312 21050 21321
rect 20994 21247 21050 21256
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20824 20058 20852 20878
rect 20916 20466 20944 20946
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 21008 19922 21036 21247
rect 21088 21140 21140 21146
rect 21088 21082 21140 21088
rect 21100 20806 21128 21082
rect 21192 20942 21220 21558
rect 21836 21146 21864 22374
rect 21824 21140 21876 21146
rect 21824 21082 21876 21088
rect 21928 21078 21956 22578
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 22020 21622 22048 21966
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 22112 21570 22140 21830
rect 22204 21690 22232 22578
rect 22296 22030 22324 22732
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 21916 21072 21968 21078
rect 21916 21014 21968 21020
rect 21180 20936 21232 20942
rect 21180 20878 21232 20884
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21088 20800 21140 20806
rect 21088 20742 21140 20748
rect 21100 20602 21128 20742
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 21468 20262 21496 20878
rect 21836 20777 21864 20878
rect 22020 20806 22048 21558
rect 22112 21542 22232 21570
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 22008 20800 22060 20806
rect 21822 20768 21878 20777
rect 22008 20742 22060 20748
rect 21822 20703 21878 20712
rect 21914 20496 21970 20505
rect 21914 20431 21970 20440
rect 21928 20262 21956 20431
rect 22112 20398 22140 20946
rect 22204 20942 22232 21542
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 22204 20806 22232 20878
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22100 20392 22152 20398
rect 22100 20334 22152 20340
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 22204 20210 22232 20742
rect 22296 20330 22324 21966
rect 22388 21026 22416 25230
rect 22480 25226 22692 25242
rect 22468 25220 22692 25226
rect 22520 25214 22692 25220
rect 22468 25162 22520 25168
rect 22756 25158 22784 26182
rect 22652 25152 22704 25158
rect 22652 25094 22704 25100
rect 22744 25152 22796 25158
rect 22744 25094 22796 25100
rect 22664 24818 22692 25094
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22664 23798 22692 24210
rect 22652 23792 22704 23798
rect 22652 23734 22704 23740
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22468 23044 22520 23050
rect 22468 22986 22520 22992
rect 22480 22642 22508 22986
rect 22468 22636 22520 22642
rect 22468 22578 22520 22584
rect 22468 21888 22520 21894
rect 22466 21856 22468 21865
rect 22520 21856 22522 21865
rect 22466 21791 22522 21800
rect 22388 20998 22508 21026
rect 22376 20936 22428 20942
rect 22374 20904 22376 20913
rect 22428 20904 22430 20913
rect 22374 20839 22430 20848
rect 22374 20360 22430 20369
rect 22284 20324 22336 20330
rect 22374 20295 22430 20304
rect 22284 20266 22336 20272
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20824 19666 20852 19722
rect 20824 19638 20944 19666
rect 20916 18970 20944 19638
rect 21928 19446 21956 20198
rect 22204 20182 22324 20210
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22098 19952 22154 19961
rect 22098 19887 22154 19896
rect 22112 19514 22140 19887
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 21916 19440 21968 19446
rect 21916 19382 21968 19388
rect 22098 19272 22154 19281
rect 22098 19207 22154 19216
rect 22112 19174 22140 19207
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20352 17264 20404 17270
rect 20352 17206 20404 17212
rect 20364 16590 20392 17206
rect 20456 16726 20484 18226
rect 20640 17610 20668 18702
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20824 17202 20852 17818
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20456 16182 20484 16662
rect 20444 16176 20496 16182
rect 20444 16118 20496 16124
rect 20548 16046 20576 17070
rect 20720 17060 20772 17066
rect 20720 17002 20772 17008
rect 20732 16726 20760 17002
rect 21008 16794 21036 18566
rect 21100 17338 21128 18906
rect 21640 18760 21692 18766
rect 22204 18714 22232 19994
rect 21640 18702 21692 18708
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 21192 17678 21220 18634
rect 21454 18048 21510 18057
rect 21454 17983 21510 17992
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20732 16250 20760 16662
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20824 16250 20852 16526
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20456 15094 20484 15846
rect 20548 15366 20576 15982
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20444 15088 20496 15094
rect 20444 15030 20496 15036
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20548 14550 20576 14758
rect 20640 14550 20668 15982
rect 20732 15910 20760 16186
rect 20916 16114 20944 16390
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 21008 16046 21036 16526
rect 20812 16040 20864 16046
rect 20812 15982 20864 15988
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20824 15026 20852 15982
rect 21100 15570 21128 17274
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20628 14544 20680 14550
rect 20628 14486 20680 14492
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20456 13938 20484 14282
rect 20548 14006 20576 14486
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20640 13954 20668 14486
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20456 13462 20484 13874
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 20548 13326 20576 13942
rect 20640 13938 20760 13954
rect 20640 13932 20772 13938
rect 20640 13926 20720 13932
rect 20720 13874 20772 13880
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20536 13184 20588 13190
rect 20456 13144 20536 13172
rect 20260 11280 20312 11286
rect 20260 11222 20312 11228
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 20088 9674 20116 11086
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 20180 10062 20208 10406
rect 20272 10266 20300 11222
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 19904 9646 20116 9674
rect 19904 9586 19932 9646
rect 20180 9586 20208 9998
rect 20272 9722 20300 10202
rect 20456 10180 20484 13144
rect 20536 13126 20588 13132
rect 20640 12646 20668 13466
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20824 12306 20852 14758
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 21100 14074 21128 14350
rect 21284 14074 21312 16186
rect 21468 16114 21496 17983
rect 21652 17882 21680 18702
rect 22112 18686 22232 18714
rect 22112 18426 22140 18686
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 22112 17678 22140 18362
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21100 13326 21128 14010
rect 21376 13954 21404 15982
rect 22020 15502 22048 16050
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 21836 14346 21864 14894
rect 22112 14482 22140 14894
rect 22204 14822 22232 18566
rect 22296 17678 22324 20182
rect 22388 19553 22416 20295
rect 22374 19544 22430 19553
rect 22374 19479 22430 19488
rect 22388 19446 22416 19479
rect 22376 19440 22428 19446
rect 22376 19382 22428 19388
rect 22374 19000 22430 19009
rect 22374 18935 22430 18944
rect 22388 18766 22416 18935
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22388 18290 22416 18702
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22296 16250 22324 16526
rect 22376 16516 22428 16522
rect 22376 16458 22428 16464
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22296 14618 22324 14758
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 22192 14068 22244 14074
rect 21284 13926 21404 13954
rect 22112 14028 22192 14056
rect 21824 13932 21876 13938
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 21192 12986 21220 13126
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 21008 12434 21036 12854
rect 20916 12406 21036 12434
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 20824 10441 20852 10474
rect 20810 10432 20866 10441
rect 20810 10367 20866 10376
rect 20536 10192 20588 10198
rect 20456 10152 20536 10180
rect 20456 10062 20484 10152
rect 20536 10134 20588 10140
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20916 9994 20944 12406
rect 21284 11898 21312 13926
rect 21824 13874 21876 13880
rect 21364 13796 21416 13802
rect 21364 13738 21416 13744
rect 21376 13326 21404 13738
rect 21836 13462 21864 13874
rect 21824 13456 21876 13462
rect 21824 13398 21876 13404
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21376 12646 21404 13262
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21560 12918 21588 13126
rect 21744 12986 21772 13262
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 21548 12912 21600 12918
rect 21548 12854 21600 12860
rect 21836 12850 21864 13398
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21468 12170 21496 12786
rect 21836 12170 21864 12786
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21824 12164 21876 12170
rect 21824 12106 21876 12112
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 22112 11778 22140 14028
rect 22192 14010 22244 14016
rect 22296 13308 22324 14418
rect 22388 13870 22416 16458
rect 22376 13864 22428 13870
rect 22480 13852 22508 20998
rect 22572 19378 22600 23258
rect 22848 22094 22876 30359
rect 22928 30252 22980 30258
rect 22928 30194 22980 30200
rect 22940 29646 22968 30194
rect 23032 29866 23060 31078
rect 23124 30569 23152 31758
rect 23110 30560 23166 30569
rect 23110 30495 23166 30504
rect 23124 30258 23152 30495
rect 23216 30326 23244 33646
rect 23308 33590 23336 35770
rect 23480 35488 23532 35494
rect 23480 35430 23532 35436
rect 23492 35290 23520 35430
rect 23480 35284 23532 35290
rect 23480 35226 23532 35232
rect 23584 35018 23612 36230
rect 23676 35834 23704 37810
rect 23768 36378 23796 37810
rect 24044 37670 24072 38150
rect 24872 38010 24900 38354
rect 25596 38276 25648 38282
rect 25596 38218 25648 38224
rect 25608 38010 25636 38218
rect 24860 38004 24912 38010
rect 24860 37946 24912 37952
rect 25596 38004 25648 38010
rect 25596 37946 25648 37952
rect 25792 37942 25820 38383
rect 26056 38354 26108 38360
rect 27620 38412 27672 38418
rect 27620 38354 27672 38360
rect 26068 38282 26096 38354
rect 29552 38344 29604 38350
rect 29552 38286 29604 38292
rect 29644 38344 29696 38350
rect 29644 38286 29696 38292
rect 26056 38276 26108 38282
rect 26056 38218 26108 38224
rect 27528 38276 27580 38282
rect 27528 38218 27580 38224
rect 29276 38276 29328 38282
rect 29276 38218 29328 38224
rect 29460 38276 29512 38282
rect 29460 38218 29512 38224
rect 26976 38208 27028 38214
rect 26976 38150 27028 38156
rect 25780 37936 25832 37942
rect 25318 37904 25374 37913
rect 25780 37878 25832 37884
rect 25318 37839 25320 37848
rect 25372 37839 25374 37848
rect 26424 37868 26476 37874
rect 25320 37810 25372 37816
rect 26424 37810 26476 37816
rect 26608 37868 26660 37874
rect 26608 37810 26660 37816
rect 25228 37800 25280 37806
rect 25228 37742 25280 37748
rect 25596 37800 25648 37806
rect 25596 37742 25648 37748
rect 26148 37800 26200 37806
rect 26148 37742 26200 37748
rect 23940 37664 23992 37670
rect 23940 37606 23992 37612
rect 24032 37664 24084 37670
rect 24032 37606 24084 37612
rect 23952 36786 23980 37606
rect 23940 36780 23992 36786
rect 23940 36722 23992 36728
rect 23940 36644 23992 36650
rect 23940 36586 23992 36592
rect 23756 36372 23808 36378
rect 23756 36314 23808 36320
rect 23952 36310 23980 36586
rect 23940 36304 23992 36310
rect 23940 36246 23992 36252
rect 23664 35828 23716 35834
rect 23664 35770 23716 35776
rect 24044 35766 24072 37606
rect 24860 37392 24912 37398
rect 25240 37369 25268 37742
rect 24860 37334 24912 37340
rect 25226 37360 25282 37369
rect 24400 37256 24452 37262
rect 24400 37198 24452 37204
rect 24124 36644 24176 36650
rect 24124 36586 24176 36592
rect 24032 35760 24084 35766
rect 24032 35702 24084 35708
rect 23756 35692 23808 35698
rect 23756 35634 23808 35640
rect 23664 35556 23716 35562
rect 23664 35498 23716 35504
rect 23676 35154 23704 35498
rect 23664 35148 23716 35154
rect 23664 35090 23716 35096
rect 23572 35012 23624 35018
rect 23572 34954 23624 34960
rect 23480 34604 23532 34610
rect 23400 34564 23480 34592
rect 23296 33584 23348 33590
rect 23296 33526 23348 33532
rect 23308 32502 23336 33526
rect 23400 32570 23428 34564
rect 23480 34546 23532 34552
rect 23478 34504 23534 34513
rect 23478 34439 23534 34448
rect 23492 33998 23520 34439
rect 23584 33998 23612 34954
rect 23768 34746 23796 35634
rect 23848 35624 23900 35630
rect 23848 35566 23900 35572
rect 23860 34950 23888 35566
rect 23940 35488 23992 35494
rect 23940 35430 23992 35436
rect 23952 35290 23980 35430
rect 23940 35284 23992 35290
rect 23940 35226 23992 35232
rect 23848 34944 23900 34950
rect 23848 34886 23900 34892
rect 23940 34944 23992 34950
rect 23940 34886 23992 34892
rect 23756 34740 23808 34746
rect 23756 34682 23808 34688
rect 23846 34640 23902 34649
rect 23676 34584 23846 34592
rect 23676 34564 23848 34584
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23572 33992 23624 33998
rect 23572 33934 23624 33940
rect 23480 33448 23532 33454
rect 23478 33416 23480 33425
rect 23532 33416 23534 33425
rect 23478 33351 23534 33360
rect 23388 32564 23440 32570
rect 23388 32506 23440 32512
rect 23296 32496 23348 32502
rect 23296 32438 23348 32444
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 23400 31958 23428 32370
rect 23388 31952 23440 31958
rect 23388 31894 23440 31900
rect 23296 31816 23348 31822
rect 23296 31758 23348 31764
rect 23308 31482 23336 31758
rect 23388 31680 23440 31686
rect 23388 31622 23440 31628
rect 23400 31521 23428 31622
rect 23386 31512 23442 31521
rect 23296 31476 23348 31482
rect 23386 31447 23442 31456
rect 23296 31418 23348 31424
rect 23296 31340 23348 31346
rect 23296 31282 23348 31288
rect 23308 30870 23336 31282
rect 23296 30864 23348 30870
rect 23296 30806 23348 30812
rect 23204 30320 23256 30326
rect 23204 30262 23256 30268
rect 23388 30320 23440 30326
rect 23388 30262 23440 30268
rect 23112 30252 23164 30258
rect 23112 30194 23164 30200
rect 23216 29866 23244 30262
rect 23400 30025 23428 30262
rect 23386 30016 23442 30025
rect 23386 29951 23442 29960
rect 23032 29838 23152 29866
rect 23216 29838 23428 29866
rect 22928 29640 22980 29646
rect 22928 29582 22980 29588
rect 23020 29164 23072 29170
rect 23020 29106 23072 29112
rect 22928 28552 22980 28558
rect 22928 28494 22980 28500
rect 22940 28014 22968 28494
rect 23032 28218 23060 29106
rect 23020 28212 23072 28218
rect 23020 28154 23072 28160
rect 22928 28008 22980 28014
rect 22928 27950 22980 27956
rect 22940 26382 22968 27950
rect 22928 26376 22980 26382
rect 22928 26318 22980 26324
rect 23124 26024 23152 29838
rect 23400 29646 23428 29838
rect 23492 29714 23520 33351
rect 23676 31906 23704 34564
rect 23900 34575 23902 34584
rect 23848 34546 23900 34552
rect 23756 34400 23808 34406
rect 23756 34342 23808 34348
rect 23768 33522 23796 34342
rect 23848 33856 23900 33862
rect 23848 33798 23900 33804
rect 23860 33522 23888 33798
rect 23756 33516 23808 33522
rect 23756 33458 23808 33464
rect 23848 33516 23900 33522
rect 23848 33458 23900 33464
rect 23952 33454 23980 34886
rect 24044 34241 24072 35702
rect 24030 34232 24086 34241
rect 24030 34167 24086 34176
rect 24044 33930 24072 34167
rect 24032 33924 24084 33930
rect 24032 33866 24084 33872
rect 23940 33448 23992 33454
rect 23940 33390 23992 33396
rect 23848 33312 23900 33318
rect 24032 33312 24084 33318
rect 23848 33254 23900 33260
rect 24030 33280 24032 33289
rect 24084 33280 24086 33289
rect 23860 32570 23888 33254
rect 24030 33215 24086 33224
rect 23940 32768 23992 32774
rect 23940 32710 23992 32716
rect 23848 32564 23900 32570
rect 23848 32506 23900 32512
rect 23952 32502 23980 32710
rect 23940 32496 23992 32502
rect 23940 32438 23992 32444
rect 24136 32434 24164 36586
rect 24308 36372 24360 36378
rect 24308 36314 24360 36320
rect 24216 33992 24268 33998
rect 24216 33934 24268 33940
rect 24124 32428 24176 32434
rect 24124 32370 24176 32376
rect 24228 32314 24256 33934
rect 24320 33153 24348 36314
rect 24306 33144 24362 33153
rect 24306 33079 24362 33088
rect 24044 32286 24256 32314
rect 23676 31878 23888 31906
rect 23572 31816 23624 31822
rect 23572 31758 23624 31764
rect 23664 31816 23716 31822
rect 23664 31758 23716 31764
rect 23584 30598 23612 31758
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23480 29708 23532 29714
rect 23480 29650 23532 29656
rect 23204 29640 23256 29646
rect 23204 29582 23256 29588
rect 23388 29640 23440 29646
rect 23676 29594 23704 31758
rect 23756 31748 23808 31754
rect 23756 31690 23808 31696
rect 23768 31113 23796 31690
rect 23754 31104 23810 31113
rect 23754 31039 23810 31048
rect 23860 30394 23888 31878
rect 23940 31816 23992 31822
rect 23940 31758 23992 31764
rect 23848 30388 23900 30394
rect 23848 30330 23900 30336
rect 23952 30054 23980 31758
rect 24044 31657 24072 32286
rect 24320 32178 24348 33079
rect 24136 32150 24348 32178
rect 24136 31890 24164 32150
rect 24412 32008 24440 37198
rect 24676 37188 24728 37194
rect 24676 37130 24728 37136
rect 24584 37120 24636 37126
rect 24584 37062 24636 37068
rect 24492 36780 24544 36786
rect 24492 36722 24544 36728
rect 24504 36310 24532 36722
rect 24596 36582 24624 37062
rect 24584 36576 24636 36582
rect 24584 36518 24636 36524
rect 24492 36304 24544 36310
rect 24492 36246 24544 36252
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 24492 33856 24544 33862
rect 24492 33798 24544 33804
rect 24504 33114 24532 33798
rect 24492 33108 24544 33114
rect 24492 33050 24544 33056
rect 24228 31980 24440 32008
rect 24124 31884 24176 31890
rect 24124 31826 24176 31832
rect 24228 31822 24256 31980
rect 24306 31920 24362 31929
rect 24596 31890 24624 36110
rect 24688 32348 24716 37130
rect 24872 35698 24900 37334
rect 25226 37295 25282 37304
rect 25136 36916 25188 36922
rect 25136 36858 25188 36864
rect 25148 36650 25176 36858
rect 25136 36644 25188 36650
rect 25136 36586 25188 36592
rect 24952 36100 25004 36106
rect 24952 36042 25004 36048
rect 24964 35698 24992 36042
rect 25148 35766 25176 36586
rect 25136 35760 25188 35766
rect 25136 35702 25188 35708
rect 24860 35692 24912 35698
rect 24860 35634 24912 35640
rect 24952 35692 25004 35698
rect 24952 35634 25004 35640
rect 25412 35692 25464 35698
rect 25412 35634 25464 35640
rect 24860 35216 24912 35222
rect 24860 35158 24912 35164
rect 24768 34400 24820 34406
rect 24768 34342 24820 34348
rect 24780 33998 24808 34342
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 24768 32360 24820 32366
rect 24688 32320 24768 32348
rect 24768 32302 24820 32308
rect 24306 31855 24362 31864
rect 24584 31884 24636 31890
rect 24320 31822 24348 31855
rect 24584 31826 24636 31832
rect 24216 31816 24268 31822
rect 24216 31758 24268 31764
rect 24308 31816 24360 31822
rect 24308 31758 24360 31764
rect 24596 31754 24624 31826
rect 24504 31726 24624 31754
rect 24030 31648 24086 31657
rect 24030 31583 24086 31592
rect 24044 31090 24072 31583
rect 24044 31062 24256 31090
rect 23940 30048 23992 30054
rect 23940 29990 23992 29996
rect 23848 29776 23900 29782
rect 23848 29718 23900 29724
rect 23388 29582 23440 29588
rect 23216 29238 23244 29582
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 23204 29232 23256 29238
rect 23204 29174 23256 29180
rect 23204 28960 23256 28966
rect 23204 28902 23256 28908
rect 23216 28082 23244 28902
rect 23308 28218 23336 29446
rect 23400 28801 23428 29582
rect 23492 29566 23704 29594
rect 23756 29640 23808 29646
rect 23756 29582 23808 29588
rect 23386 28792 23442 28801
rect 23386 28727 23442 28736
rect 23296 28212 23348 28218
rect 23296 28154 23348 28160
rect 23204 28076 23256 28082
rect 23204 28018 23256 28024
rect 23388 28076 23440 28082
rect 23388 28018 23440 28024
rect 23400 27674 23428 28018
rect 23388 27668 23440 27674
rect 23388 27610 23440 27616
rect 23492 27062 23520 29566
rect 23572 29504 23624 29510
rect 23572 29446 23624 29452
rect 23584 29073 23612 29446
rect 23676 29238 23704 29566
rect 23664 29232 23716 29238
rect 23664 29174 23716 29180
rect 23570 29064 23626 29073
rect 23570 28999 23626 29008
rect 23768 28558 23796 29582
rect 23860 29306 23888 29718
rect 23848 29300 23900 29306
rect 23848 29242 23900 29248
rect 23952 29170 23980 29990
rect 24124 29844 24176 29850
rect 24124 29786 24176 29792
rect 23940 29164 23992 29170
rect 23940 29106 23992 29112
rect 23940 29028 23992 29034
rect 23940 28970 23992 28976
rect 23756 28552 23808 28558
rect 23756 28494 23808 28500
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23768 28082 23796 28358
rect 23572 28076 23624 28082
rect 23572 28018 23624 28024
rect 23756 28076 23808 28082
rect 23756 28018 23808 28024
rect 23584 27606 23612 28018
rect 23572 27600 23624 27606
rect 23572 27542 23624 27548
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23480 27056 23532 27062
rect 23480 26998 23532 27004
rect 23296 26376 23348 26382
rect 23296 26318 23348 26324
rect 23124 25996 23244 26024
rect 23020 25968 23072 25974
rect 23020 25910 23072 25916
rect 23110 25936 23166 25945
rect 22928 25832 22980 25838
rect 22928 25774 22980 25780
rect 22940 24954 22968 25774
rect 23032 24954 23060 25910
rect 23110 25871 23112 25880
rect 23164 25871 23166 25880
rect 23112 25842 23164 25848
rect 23112 25696 23164 25702
rect 23112 25638 23164 25644
rect 23124 25362 23152 25638
rect 23112 25356 23164 25362
rect 23112 25298 23164 25304
rect 22928 24948 22980 24954
rect 22928 24890 22980 24896
rect 23020 24948 23072 24954
rect 23020 24890 23072 24896
rect 23112 23860 23164 23866
rect 23112 23802 23164 23808
rect 22928 23724 22980 23730
rect 22928 23666 22980 23672
rect 23020 23724 23072 23730
rect 23020 23666 23072 23672
rect 22940 23118 22968 23666
rect 23032 23118 23060 23666
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 23020 23112 23072 23118
rect 23020 23054 23072 23060
rect 22940 22778 22968 23054
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 22756 22066 22876 22094
rect 22650 21720 22706 21729
rect 22650 21655 22706 21664
rect 22664 19854 22692 21655
rect 22652 19848 22704 19854
rect 22652 19790 22704 19796
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22572 18290 22600 19314
rect 22652 18964 22704 18970
rect 22652 18906 22704 18912
rect 22664 18358 22692 18906
rect 22652 18352 22704 18358
rect 22652 18294 22704 18300
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22650 17912 22706 17921
rect 22756 17882 22784 22066
rect 23032 21962 23060 23054
rect 23020 21956 23072 21962
rect 23020 21898 23072 21904
rect 22834 21448 22890 21457
rect 23124 21434 23152 23802
rect 22834 21383 22890 21392
rect 22928 21412 22980 21418
rect 22848 20806 22876 21383
rect 22928 21354 22980 21360
rect 23032 21406 23152 21434
rect 22940 21321 22968 21354
rect 22926 21312 22982 21321
rect 22926 21247 22982 21256
rect 22928 21004 22980 21010
rect 22928 20946 22980 20952
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22940 20058 22968 20946
rect 22928 20052 22980 20058
rect 22928 19994 22980 20000
rect 22836 19780 22888 19786
rect 22836 19722 22888 19728
rect 22848 19514 22876 19722
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22650 17847 22706 17856
rect 22744 17876 22796 17882
rect 22664 15570 22692 17847
rect 22744 17818 22796 17824
rect 22928 17196 22980 17202
rect 22928 17138 22980 17144
rect 22940 16590 22968 17138
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 22836 16516 22888 16522
rect 22836 16458 22888 16464
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22560 13864 22612 13870
rect 22480 13824 22560 13852
rect 22376 13806 22428 13812
rect 22560 13806 22612 13812
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22376 13320 22428 13326
rect 22296 13280 22376 13308
rect 22376 13262 22428 13268
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22204 12782 22232 13126
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22204 11898 22232 12718
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22296 11830 22324 12718
rect 22388 12442 22416 13262
rect 22572 12714 22600 13670
rect 22560 12708 22612 12714
rect 22560 12650 22612 12656
rect 22376 12436 22428 12442
rect 22664 12434 22692 15506
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22756 13870 22784 14486
rect 22848 14414 22876 16458
rect 23032 16182 23060 21406
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23124 21078 23152 21286
rect 23112 21072 23164 21078
rect 23112 21014 23164 21020
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 23124 17134 23152 19314
rect 23216 18970 23244 25996
rect 23308 23322 23336 26318
rect 23388 26240 23440 26246
rect 23388 26182 23440 26188
rect 23400 23866 23428 26182
rect 23478 25528 23534 25537
rect 23584 25498 23612 27406
rect 23756 26240 23808 26246
rect 23756 26182 23808 26188
rect 23768 26042 23796 26182
rect 23756 26036 23808 26042
rect 23756 25978 23808 25984
rect 23952 25838 23980 28970
rect 24032 28960 24084 28966
rect 24032 28902 24084 28908
rect 24044 28082 24072 28902
rect 24032 28076 24084 28082
rect 24032 28018 24084 28024
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23940 25832 23992 25838
rect 23940 25774 23992 25780
rect 23478 25463 23534 25472
rect 23572 25492 23624 25498
rect 23492 25362 23520 25463
rect 23572 25434 23624 25440
rect 23480 25356 23532 25362
rect 23532 25316 23612 25344
rect 23480 25298 23532 25304
rect 23584 24818 23612 25316
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23572 24812 23624 24818
rect 23572 24754 23624 24760
rect 23492 24206 23520 24754
rect 23676 24410 23704 25774
rect 23848 24744 23900 24750
rect 23848 24686 23900 24692
rect 23664 24404 23716 24410
rect 23664 24346 23716 24352
rect 23572 24336 23624 24342
rect 23572 24278 23624 24284
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23400 22642 23428 23258
rect 23492 23254 23520 24142
rect 23480 23248 23532 23254
rect 23480 23190 23532 23196
rect 23584 22642 23612 24278
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23768 23730 23796 24142
rect 23860 23730 23888 24686
rect 23952 24449 23980 25774
rect 24136 25702 24164 29786
rect 24228 28937 24256 31062
rect 24400 30932 24452 30938
rect 24400 30874 24452 30880
rect 24412 29850 24440 30874
rect 24400 29844 24452 29850
rect 24400 29786 24452 29792
rect 24308 29640 24360 29646
rect 24308 29582 24360 29588
rect 24214 28928 24270 28937
rect 24214 28863 24270 28872
rect 24228 28218 24256 28863
rect 24216 28212 24268 28218
rect 24216 28154 24268 28160
rect 24216 27872 24268 27878
rect 24216 27814 24268 27820
rect 24228 27674 24256 27814
rect 24216 27668 24268 27674
rect 24216 27610 24268 27616
rect 24320 25906 24348 29582
rect 24504 28626 24532 31726
rect 24780 31686 24808 32302
rect 24768 31680 24820 31686
rect 24768 31622 24820 31628
rect 24584 31272 24636 31278
rect 24584 31214 24636 31220
rect 24596 30802 24624 31214
rect 24584 30796 24636 30802
rect 24584 30738 24636 30744
rect 24584 30660 24636 30666
rect 24584 30602 24636 30608
rect 24596 29714 24624 30602
rect 24676 30320 24728 30326
rect 24676 30262 24728 30268
rect 24688 29714 24716 30262
rect 24584 29708 24636 29714
rect 24584 29650 24636 29656
rect 24676 29708 24728 29714
rect 24676 29650 24728 29656
rect 24492 28620 24544 28626
rect 24492 28562 24544 28568
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24400 28416 24452 28422
rect 24400 28358 24452 28364
rect 24412 28082 24440 28358
rect 24688 28082 24716 28494
rect 24780 28490 24808 31622
rect 24768 28484 24820 28490
rect 24768 28426 24820 28432
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24676 28076 24728 28082
rect 24676 28018 24728 28024
rect 24492 27872 24544 27878
rect 24398 27840 24454 27849
rect 24492 27814 24544 27820
rect 24398 27775 24454 27784
rect 24412 27674 24440 27775
rect 24400 27668 24452 27674
rect 24400 27610 24452 27616
rect 24504 26382 24532 27814
rect 24780 27130 24808 28426
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 24676 26988 24728 26994
rect 24596 26948 24676 26976
rect 24492 26376 24544 26382
rect 24492 26318 24544 26324
rect 24596 26194 24624 26948
rect 24676 26930 24728 26936
rect 24768 26920 24820 26926
rect 24768 26862 24820 26868
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24504 26166 24624 26194
rect 24308 25900 24360 25906
rect 24308 25842 24360 25848
rect 24216 25832 24268 25838
rect 24216 25774 24268 25780
rect 24124 25696 24176 25702
rect 24124 25638 24176 25644
rect 24228 25430 24256 25774
rect 24320 25673 24348 25842
rect 24306 25664 24362 25673
rect 24306 25599 24362 25608
rect 24216 25424 24268 25430
rect 24216 25366 24268 25372
rect 24216 24676 24268 24682
rect 24216 24618 24268 24624
rect 23938 24440 23994 24449
rect 23938 24375 23994 24384
rect 24228 24206 24256 24618
rect 23940 24200 23992 24206
rect 23940 24142 23992 24148
rect 24216 24200 24268 24206
rect 24216 24142 24268 24148
rect 23756 23724 23808 23730
rect 23756 23666 23808 23672
rect 23848 23724 23900 23730
rect 23848 23666 23900 23672
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23676 22778 23704 22918
rect 23768 22778 23796 23666
rect 23860 23186 23888 23666
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23756 22772 23808 22778
rect 23756 22714 23808 22720
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 23308 21486 23336 22578
rect 23584 22166 23612 22578
rect 23572 22160 23624 22166
rect 23572 22102 23624 22108
rect 23480 22024 23532 22030
rect 23480 21966 23532 21972
rect 23388 21956 23440 21962
rect 23388 21898 23440 21904
rect 23296 21480 23348 21486
rect 23296 21422 23348 21428
rect 23308 20602 23336 21422
rect 23400 21010 23428 21898
rect 23492 21418 23520 21966
rect 23860 21622 23888 23122
rect 23952 22506 23980 24142
rect 24400 23656 24452 23662
rect 24306 23624 24362 23633
rect 24400 23598 24452 23604
rect 24306 23559 24308 23568
rect 24360 23559 24362 23568
rect 24308 23530 24360 23536
rect 24412 23118 24440 23598
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 24400 23112 24452 23118
rect 24400 23054 24452 23060
rect 24044 22642 24072 23054
rect 24124 23044 24176 23050
rect 24124 22986 24176 22992
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 23940 22500 23992 22506
rect 23940 22442 23992 22448
rect 24044 22098 24072 22578
rect 24136 22574 24164 22986
rect 24124 22568 24176 22574
rect 24124 22510 24176 22516
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 24504 22030 24532 26166
rect 24688 25906 24716 26318
rect 24780 26042 24808 26862
rect 24768 26036 24820 26042
rect 24768 25978 24820 25984
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24768 25900 24820 25906
rect 24768 25842 24820 25848
rect 24688 24342 24716 25842
rect 24780 25498 24808 25842
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24676 24336 24728 24342
rect 24676 24278 24728 24284
rect 24688 23712 24716 24278
rect 24768 23724 24820 23730
rect 24688 23684 24768 23712
rect 24768 23666 24820 23672
rect 24872 23186 24900 35158
rect 24964 34474 24992 35634
rect 25424 35290 25452 35634
rect 25504 35488 25556 35494
rect 25504 35430 25556 35436
rect 25412 35284 25464 35290
rect 25412 35226 25464 35232
rect 25320 35080 25372 35086
rect 25320 35022 25372 35028
rect 25228 34944 25280 34950
rect 25228 34886 25280 34892
rect 24952 34468 25004 34474
rect 24952 34410 25004 34416
rect 24964 31686 24992 34410
rect 25136 32020 25188 32026
rect 25056 31980 25136 32008
rect 25056 31822 25084 31980
rect 25136 31962 25188 31968
rect 25044 31816 25096 31822
rect 25044 31758 25096 31764
rect 25136 31816 25188 31822
rect 25136 31758 25188 31764
rect 24952 31680 25004 31686
rect 24952 31622 25004 31628
rect 25148 30938 25176 31758
rect 25136 30932 25188 30938
rect 25136 30874 25188 30880
rect 25134 30560 25190 30569
rect 25134 30495 25190 30504
rect 24950 29880 25006 29889
rect 24950 29815 25006 29824
rect 24964 29646 24992 29815
rect 25148 29782 25176 30495
rect 25136 29776 25188 29782
rect 25136 29718 25188 29724
rect 24952 29640 25004 29646
rect 24952 29582 25004 29588
rect 24952 28552 25004 28558
rect 24952 28494 25004 28500
rect 24964 28422 24992 28494
rect 24952 28416 25004 28422
rect 24952 28358 25004 28364
rect 25134 26072 25190 26081
rect 25056 26016 25134 26024
rect 25056 25996 25136 26016
rect 24950 25800 25006 25809
rect 24950 25735 24952 25744
rect 25004 25735 25006 25744
rect 24952 25706 25004 25712
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24858 22672 24914 22681
rect 24858 22607 24914 22616
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24584 22160 24636 22166
rect 24584 22102 24636 22108
rect 24674 22128 24730 22137
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 23848 21616 23900 21622
rect 23848 21558 23900 21564
rect 23480 21412 23532 21418
rect 23480 21354 23532 21360
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23400 20233 23428 20538
rect 24412 20466 24440 20878
rect 24504 20874 24532 21966
rect 24492 20868 24544 20874
rect 24492 20810 24544 20816
rect 24596 20466 24624 22102
rect 24674 22063 24730 22072
rect 24688 21690 24716 22063
rect 24780 22030 24808 22374
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24872 21729 24900 22607
rect 24952 22160 25004 22166
rect 24952 22102 25004 22108
rect 24858 21720 24914 21729
rect 24676 21684 24728 21690
rect 24858 21655 24914 21664
rect 24676 21626 24728 21632
rect 24768 21616 24820 21622
rect 24768 21558 24820 21564
rect 24400 20460 24452 20466
rect 24584 20460 24636 20466
rect 24400 20402 24452 20408
rect 24504 20420 24584 20448
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23386 20224 23442 20233
rect 23386 20159 23442 20168
rect 23400 20058 23428 20159
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23584 19854 23612 20334
rect 24032 20256 24084 20262
rect 24032 20198 24084 20204
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23940 19916 23992 19922
rect 23940 19858 23992 19864
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23388 19848 23440 19854
rect 23572 19848 23624 19854
rect 23388 19790 23440 19796
rect 23478 19816 23534 19825
rect 23204 18964 23256 18970
rect 23204 18906 23256 18912
rect 23308 17882 23336 19790
rect 23400 19689 23428 19790
rect 23572 19790 23624 19796
rect 23478 19751 23534 19760
rect 23492 19718 23520 19751
rect 23480 19712 23532 19718
rect 23386 19680 23442 19689
rect 23480 19654 23532 19660
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23386 19615 23442 19624
rect 23400 19378 23428 19615
rect 23480 19440 23532 19446
rect 23480 19382 23532 19388
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23492 18834 23520 19382
rect 23584 18873 23612 19654
rect 23860 19514 23888 19858
rect 23952 19514 23980 19858
rect 24044 19825 24072 20198
rect 24136 20058 24164 20198
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24504 19854 24532 20420
rect 24584 20402 24636 20408
rect 24676 20324 24728 20330
rect 24676 20266 24728 20272
rect 24688 19854 24716 20266
rect 24780 19854 24808 21558
rect 24858 21176 24914 21185
rect 24858 21111 24914 21120
rect 24872 20942 24900 21111
rect 24964 21010 24992 22102
rect 25056 21434 25084 25996
rect 25188 26007 25190 26016
rect 25136 25978 25188 25984
rect 25136 25900 25188 25906
rect 25136 25842 25188 25848
rect 25148 25537 25176 25842
rect 25134 25528 25190 25537
rect 25134 25463 25190 25472
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 25148 23730 25176 24754
rect 25136 23724 25188 23730
rect 25136 23666 25188 23672
rect 25148 23118 25176 23666
rect 25136 23112 25188 23118
rect 25136 23054 25188 23060
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25148 21554 25176 21626
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25056 21406 25176 21434
rect 25042 21176 25098 21185
rect 25042 21111 25044 21120
rect 25096 21111 25098 21120
rect 25044 21082 25096 21088
rect 25148 21026 25176 21406
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 25056 20998 25176 21026
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24872 20466 24900 20742
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 24492 19848 24544 19854
rect 24030 19816 24086 19825
rect 24492 19790 24544 19796
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24030 19751 24086 19760
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 23570 18864 23626 18873
rect 23480 18828 23532 18834
rect 23570 18799 23626 18808
rect 23480 18770 23532 18776
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23386 17912 23442 17921
rect 23296 17876 23348 17882
rect 23386 17847 23442 17856
rect 23296 17818 23348 17824
rect 23202 17640 23258 17649
rect 23202 17575 23258 17584
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 23216 16658 23244 17575
rect 23308 17338 23336 17818
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 23296 17060 23348 17066
rect 23296 17002 23348 17008
rect 23204 16652 23256 16658
rect 23204 16594 23256 16600
rect 23308 16561 23336 17002
rect 23400 16590 23428 17847
rect 23676 17814 23704 18158
rect 23664 17808 23716 17814
rect 23664 17750 23716 17756
rect 23480 17740 23532 17746
rect 23480 17682 23532 17688
rect 23492 17338 23520 17682
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23388 16584 23440 16590
rect 23294 16552 23350 16561
rect 23204 16516 23256 16522
rect 23388 16526 23440 16532
rect 23294 16487 23296 16496
rect 23204 16458 23256 16464
rect 23348 16487 23350 16496
rect 23756 16516 23808 16522
rect 23296 16458 23348 16464
rect 23756 16458 23808 16464
rect 23020 16176 23072 16182
rect 23020 16118 23072 16124
rect 23032 15502 23060 16118
rect 23216 16114 23244 16458
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 23216 15706 23244 16050
rect 23768 16017 23796 16458
rect 23754 16008 23810 16017
rect 23754 15943 23810 15952
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 23952 15502 23980 18226
rect 24044 17678 24072 19751
rect 24504 19446 24532 19790
rect 24860 19780 24912 19786
rect 24860 19722 24912 19728
rect 24768 19508 24820 19514
rect 24872 19496 24900 19722
rect 24820 19468 24900 19496
rect 24768 19450 24820 19456
rect 24492 19440 24544 19446
rect 24492 19382 24544 19388
rect 24308 19304 24360 19310
rect 24306 19272 24308 19281
rect 24360 19272 24362 19281
rect 24306 19207 24362 19216
rect 24124 19168 24176 19174
rect 24124 19110 24176 19116
rect 24032 17672 24084 17678
rect 24032 17614 24084 17620
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 23202 15056 23258 15065
rect 23202 14991 23204 15000
rect 23256 14991 23258 15000
rect 23204 14962 23256 14968
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22848 14074 22876 14214
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 22744 13864 22796 13870
rect 22796 13824 22876 13852
rect 22744 13806 22796 13812
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22756 13462 22784 13670
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22376 12378 22428 12384
rect 22572 12406 22692 12434
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22284 11824 22336 11830
rect 21836 11286 21864 11766
rect 22112 11750 22232 11778
rect 22284 11766 22336 11772
rect 22100 11620 22152 11626
rect 22100 11562 22152 11568
rect 21824 11280 21876 11286
rect 21824 11222 21876 11228
rect 22112 11082 22140 11562
rect 20996 11076 21048 11082
rect 20996 11018 21048 11024
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 21008 10742 21036 11018
rect 21456 11008 21508 11014
rect 21454 10976 21456 10985
rect 21824 11008 21876 11014
rect 21508 10976 21510 10985
rect 21824 10950 21876 10956
rect 21454 10911 21510 10920
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 20996 10736 21048 10742
rect 21560 10713 21588 10746
rect 21546 10704 21602 10713
rect 20996 10678 21048 10684
rect 21100 10662 21312 10690
rect 21100 10470 21128 10662
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 21284 10554 21312 10662
rect 21836 10690 21864 10950
rect 21546 10639 21602 10648
rect 21652 10662 21864 10690
rect 21652 10606 21680 10662
rect 21640 10600 21692 10606
rect 21284 10548 21640 10554
rect 21284 10542 21692 10548
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 20352 9988 20404 9994
rect 20352 9930 20404 9936
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20364 9897 20392 9930
rect 20350 9888 20406 9897
rect 20350 9823 20406 9832
rect 20260 9716 20312 9722
rect 20312 9664 20392 9674
rect 20260 9658 20392 9664
rect 20272 9646 20392 9658
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 19076 9178 19104 9386
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 18984 8634 19012 9046
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18970 8528 19026 8537
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18880 8492 18932 8498
rect 18970 8463 18972 8472
rect 18880 8434 18932 8440
rect 19024 8463 19026 8472
rect 18972 8434 19024 8440
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17328 6934 17356 7686
rect 17788 7410 17816 7822
rect 18616 7546 18644 8434
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17788 7002 17816 7346
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17316 6928 17368 6934
rect 17316 6870 17368 6876
rect 17880 6866 17908 7142
rect 18064 7002 18092 7142
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18234 6896 18290 6905
rect 17868 6860 17920 6866
rect 18234 6831 18290 6840
rect 17868 6802 17920 6808
rect 17880 6458 17908 6802
rect 18248 6798 18276 6831
rect 18616 6798 18644 7482
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18708 7342 18736 7414
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 18248 6338 18276 6734
rect 18616 6390 18644 6734
rect 18708 6458 18736 7278
rect 18984 6798 19012 8434
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18156 6322 18276 6338
rect 18604 6384 18656 6390
rect 18604 6326 18656 6332
rect 18984 6322 19012 6734
rect 19352 6458 19380 9318
rect 19444 8090 19472 9454
rect 19904 9058 19932 9522
rect 20260 9512 20312 9518
rect 20260 9454 20312 9460
rect 19904 9030 20208 9058
rect 20272 9042 20300 9454
rect 20364 9042 20392 9646
rect 19904 8974 19932 9030
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19996 8498 20024 8910
rect 20180 8906 20208 9030
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20076 8900 20128 8906
rect 20076 8842 20128 8848
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19536 7954 19564 8230
rect 19524 7948 19576 7954
rect 19444 7908 19524 7936
rect 19444 7342 19472 7908
rect 19524 7890 19576 7896
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6458 20024 6802
rect 20088 6458 20116 8842
rect 20180 8430 20208 8842
rect 20272 8634 20300 8978
rect 20640 8974 20668 9930
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 18144 6316 18276 6322
rect 18196 6310 18276 6316
rect 18972 6316 19024 6322
rect 18144 6258 18196 6264
rect 18972 6258 19024 6264
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 18156 5914 18184 6122
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 19536 5778 19564 6054
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19352 5302 19380 5714
rect 19536 5658 19564 5714
rect 19444 5630 19564 5658
rect 19720 5642 19748 6258
rect 20088 5914 20116 6394
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 19708 5636 19760 5642
rect 19444 5302 19472 5630
rect 19708 5578 19760 5584
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19996 4826 20024 5510
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 20088 4554 20116 5646
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20180 4826 20208 5306
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20272 4690 20300 7958
rect 20260 4684 20312 4690
rect 20260 4626 20312 4632
rect 20364 4622 20392 8774
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20548 7206 20576 7686
rect 20640 7410 20668 7890
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 20548 5710 20576 7142
rect 20640 6798 20668 7346
rect 20916 7206 20944 9930
rect 21100 9178 21128 10406
rect 21192 10062 21220 10542
rect 21284 10526 21680 10542
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21652 10062 21680 10406
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21640 10056 21692 10062
rect 21744 10044 21772 10662
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 21824 10532 21876 10538
rect 21824 10474 21876 10480
rect 21836 10266 21864 10474
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21824 10056 21876 10062
rect 21744 10016 21824 10044
rect 21640 9998 21692 10004
rect 21824 9998 21876 10004
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21100 7342 21128 9114
rect 21652 8566 21680 9998
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21836 8634 21864 8774
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 21652 7886 21680 8502
rect 21836 7886 21864 8570
rect 21928 8362 21956 10542
rect 22204 10062 22232 11750
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22296 10062 22324 11222
rect 22388 11218 22416 12038
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22572 10985 22600 12406
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22558 10976 22614 10985
rect 22558 10911 22614 10920
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22388 10470 22416 10610
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22480 10266 22508 10610
rect 22376 10260 22428 10266
rect 22376 10202 22428 10208
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22192 10056 22244 10062
rect 22192 9998 22244 10004
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21916 8356 21968 8362
rect 21916 8298 21968 8304
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21088 7336 21140 7342
rect 21088 7278 21140 7284
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 21100 6882 21128 7278
rect 21284 7002 21312 7278
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21100 6854 21312 6882
rect 21284 6798 21312 6854
rect 21376 6798 21404 7482
rect 22020 7274 22048 8434
rect 22112 7750 22140 9114
rect 22204 9042 22232 9998
rect 22388 9722 22416 10202
rect 22572 10062 22600 10911
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22282 9616 22338 9625
rect 22282 9551 22338 9560
rect 22296 9450 22324 9551
rect 22284 9444 22336 9450
rect 22284 9386 22336 9392
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 22572 8974 22600 9318
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22284 8900 22336 8906
rect 22284 8842 22336 8848
rect 22296 7954 22324 8842
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22388 7954 22416 8230
rect 22664 8106 22692 11834
rect 22848 10674 22876 13824
rect 22928 13796 22980 13802
rect 22980 13756 23060 13784
rect 22928 13738 22980 13744
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 22940 10742 22968 13398
rect 23032 12306 23060 13756
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23032 12170 23060 12242
rect 23020 12164 23072 12170
rect 23020 12106 23072 12112
rect 22928 10736 22980 10742
rect 23032 10724 23060 12106
rect 23124 11218 23152 14554
rect 23216 14482 23244 14962
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 23216 14006 23244 14282
rect 23204 14000 23256 14006
rect 23204 13942 23256 13948
rect 23216 13870 23244 13942
rect 23492 13870 23520 14350
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23664 13864 23716 13870
rect 23848 13864 23900 13870
rect 23716 13824 23796 13852
rect 23664 13806 23716 13812
rect 23216 13410 23244 13806
rect 23216 13382 23336 13410
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23216 12850 23244 13262
rect 23204 12844 23256 12850
rect 23204 12786 23256 12792
rect 23216 12238 23244 12786
rect 23308 12306 23336 13382
rect 23572 12436 23624 12442
rect 23572 12378 23624 12384
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23112 11212 23164 11218
rect 23112 11154 23164 11160
rect 23308 11082 23336 12242
rect 23584 11762 23612 12378
rect 23572 11756 23624 11762
rect 23624 11716 23704 11744
rect 23572 11698 23624 11704
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 23492 11558 23520 11630
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 23112 10736 23164 10742
rect 23032 10713 23112 10724
rect 22928 10678 22980 10684
rect 23018 10704 23112 10713
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22756 10266 22784 10406
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 22940 9926 22968 10678
rect 23074 10696 23112 10704
rect 23112 10678 23164 10684
rect 23018 10639 23074 10648
rect 23308 10606 23336 11018
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23400 10742 23428 10950
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 23296 10600 23348 10606
rect 23296 10542 23348 10548
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22744 9444 22796 9450
rect 22744 9386 22796 9392
rect 22480 8078 22692 8106
rect 22284 7948 22336 7954
rect 22284 7890 22336 7896
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22376 7812 22428 7818
rect 22376 7754 22428 7760
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22296 7546 22324 7686
rect 22388 7546 22416 7754
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22480 7426 22508 8078
rect 22756 8022 22784 9386
rect 22940 9110 22968 9862
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 22928 9104 22980 9110
rect 22834 9072 22890 9081
rect 22928 9046 22980 9052
rect 22834 9007 22890 9016
rect 22652 8016 22704 8022
rect 22652 7958 22704 7964
rect 22744 8016 22796 8022
rect 22744 7958 22796 7964
rect 22664 7886 22692 7958
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22560 7812 22612 7818
rect 22560 7754 22612 7760
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22192 7404 22244 7410
rect 22296 7398 22508 7426
rect 22296 7392 22324 7398
rect 22244 7364 22324 7392
rect 22192 7346 22244 7352
rect 22008 7268 22060 7274
rect 22008 7210 22060 7216
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 22112 6730 22140 7346
rect 22480 7002 22508 7398
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20456 5370 20484 5646
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20548 4554 20576 5646
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 21008 5302 21036 5510
rect 20996 5296 21048 5302
rect 20996 5238 21048 5244
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 20916 4826 20944 5170
rect 21008 4826 21036 5238
rect 22388 5166 22416 6598
rect 22572 6390 22600 7754
rect 22560 6384 22612 6390
rect 22560 6326 22612 6332
rect 22664 6322 22692 7822
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22664 5710 22692 6258
rect 22848 5914 22876 9007
rect 23032 8974 23060 9658
rect 23124 9110 23152 10542
rect 23400 9586 23428 10678
rect 23492 10674 23520 11290
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23492 9722 23520 10610
rect 23584 9722 23612 11222
rect 23676 11150 23704 11716
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23768 10606 23796 13824
rect 23848 13806 23900 13812
rect 23860 13462 23888 13806
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 23480 9716 23532 9722
rect 23480 9658 23532 9664
rect 23572 9716 23624 9722
rect 23572 9658 23624 9664
rect 23756 9648 23808 9654
rect 23756 9590 23808 9596
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23296 9512 23348 9518
rect 23296 9454 23348 9460
rect 23112 9104 23164 9110
rect 23112 9046 23164 9052
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 23124 8378 23152 9046
rect 23308 8906 23336 9454
rect 23400 8974 23428 9522
rect 23768 9353 23796 9590
rect 23754 9344 23810 9353
rect 23754 9279 23810 9288
rect 23768 8974 23796 9279
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23756 8968 23808 8974
rect 23756 8910 23808 8916
rect 23296 8900 23348 8906
rect 23296 8842 23348 8848
rect 23572 8832 23624 8838
rect 23572 8774 23624 8780
rect 23584 8634 23612 8774
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23860 8498 23888 12174
rect 23952 11694 23980 15438
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23952 9217 23980 11630
rect 24044 10470 24072 17614
rect 24136 14890 24164 19110
rect 24676 18148 24728 18154
rect 24676 18090 24728 18096
rect 24688 17746 24716 18090
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24688 17105 24716 17682
rect 24780 17678 24808 19450
rect 24964 19145 24992 20198
rect 24950 19136 25006 19145
rect 24950 19071 25006 19080
rect 25056 18290 25084 20998
rect 25240 20466 25268 34886
rect 25332 34746 25360 35022
rect 25320 34740 25372 34746
rect 25320 34682 25372 34688
rect 25332 33590 25360 34682
rect 25424 33998 25452 35226
rect 25516 35086 25544 35430
rect 25504 35080 25556 35086
rect 25504 35022 25556 35028
rect 25608 34950 25636 37742
rect 25688 37664 25740 37670
rect 25688 37606 25740 37612
rect 25596 34944 25648 34950
rect 25596 34886 25648 34892
rect 25412 33992 25464 33998
rect 25412 33934 25464 33940
rect 25412 33856 25464 33862
rect 25412 33798 25464 33804
rect 25320 33584 25372 33590
rect 25320 33526 25372 33532
rect 25332 32314 25360 33526
rect 25424 33454 25452 33798
rect 25412 33448 25464 33454
rect 25412 33390 25464 33396
rect 25412 33312 25464 33318
rect 25410 33280 25412 33289
rect 25464 33280 25466 33289
rect 25410 33215 25466 33224
rect 25332 32286 25452 32314
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25332 31822 25360 32166
rect 25320 31816 25372 31822
rect 25320 31758 25372 31764
rect 25424 31346 25452 32286
rect 25504 31952 25556 31958
rect 25504 31894 25556 31900
rect 25516 31793 25544 31894
rect 25502 31784 25558 31793
rect 25502 31719 25558 31728
rect 25596 31680 25648 31686
rect 25596 31622 25648 31628
rect 25504 31408 25556 31414
rect 25504 31350 25556 31356
rect 25412 31340 25464 31346
rect 25412 31282 25464 31288
rect 25424 31142 25452 31282
rect 25412 31136 25464 31142
rect 25412 31078 25464 31084
rect 25412 30728 25464 30734
rect 25412 30670 25464 30676
rect 25320 30048 25372 30054
rect 25320 29990 25372 29996
rect 25332 28558 25360 29990
rect 25424 29170 25452 30670
rect 25412 29164 25464 29170
rect 25412 29106 25464 29112
rect 25412 28960 25464 28966
rect 25412 28902 25464 28908
rect 25320 28552 25372 28558
rect 25320 28494 25372 28500
rect 25424 26976 25452 28902
rect 25516 27606 25544 31350
rect 25608 31346 25636 31622
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25596 29164 25648 29170
rect 25596 29106 25648 29112
rect 25608 28762 25636 29106
rect 25596 28756 25648 28762
rect 25596 28698 25648 28704
rect 25596 28552 25648 28558
rect 25596 28494 25648 28500
rect 25504 27600 25556 27606
rect 25504 27542 25556 27548
rect 25608 27452 25636 28494
rect 25332 26948 25452 26976
rect 25516 27424 25636 27452
rect 25332 26382 25360 26948
rect 25410 26888 25466 26897
rect 25410 26823 25466 26832
rect 25424 26586 25452 26823
rect 25516 26586 25544 27424
rect 25412 26580 25464 26586
rect 25412 26522 25464 26528
rect 25504 26580 25556 26586
rect 25504 26522 25556 26528
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25332 26042 25360 26318
rect 25320 26036 25372 26042
rect 25320 25978 25372 25984
rect 25516 25906 25544 26522
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25504 25900 25556 25906
rect 25504 25842 25556 25848
rect 25412 25832 25464 25838
rect 25412 25774 25464 25780
rect 25320 25696 25372 25702
rect 25320 25638 25372 25644
rect 25332 25158 25360 25638
rect 25320 25152 25372 25158
rect 25320 25094 25372 25100
rect 25424 24886 25452 25774
rect 25608 25770 25636 26318
rect 25596 25764 25648 25770
rect 25596 25706 25648 25712
rect 25700 25514 25728 37606
rect 25964 36168 26016 36174
rect 25964 36110 26016 36116
rect 25976 35834 26004 36110
rect 26056 36032 26108 36038
rect 26056 35974 26108 35980
rect 26068 35834 26096 35974
rect 25964 35828 26016 35834
rect 25964 35770 26016 35776
rect 26056 35828 26108 35834
rect 26056 35770 26108 35776
rect 25872 35692 25924 35698
rect 25872 35634 25924 35640
rect 25884 35562 25912 35634
rect 25872 35556 25924 35562
rect 25872 35498 25924 35504
rect 25976 34678 26004 35770
rect 26056 35692 26108 35698
rect 26056 35634 26108 35640
rect 25964 34672 26016 34678
rect 25964 34614 26016 34620
rect 25964 33992 26016 33998
rect 26068 33980 26096 35634
rect 26160 35222 26188 37742
rect 26436 37466 26464 37810
rect 26620 37466 26648 37810
rect 26424 37460 26476 37466
rect 26424 37402 26476 37408
rect 26608 37460 26660 37466
rect 26608 37402 26660 37408
rect 26988 37194 27016 38150
rect 27540 38010 27568 38218
rect 28540 38208 28592 38214
rect 28540 38150 28592 38156
rect 27528 38004 27580 38010
rect 27528 37946 27580 37952
rect 27068 37800 27120 37806
rect 27068 37742 27120 37748
rect 27988 37800 28040 37806
rect 27988 37742 28040 37748
rect 26976 37188 27028 37194
rect 26976 37130 27028 37136
rect 26240 36576 26292 36582
rect 26240 36518 26292 36524
rect 26148 35216 26200 35222
rect 26148 35158 26200 35164
rect 26148 34672 26200 34678
rect 26148 34614 26200 34620
rect 26160 33998 26188 34614
rect 26016 33952 26096 33980
rect 26148 33992 26200 33998
rect 25964 33934 26016 33940
rect 26148 33934 26200 33940
rect 25976 32434 26004 33934
rect 26160 33046 26188 33934
rect 26148 33040 26200 33046
rect 26148 32982 26200 32988
rect 25964 32428 26016 32434
rect 25964 32370 26016 32376
rect 25780 32360 25832 32366
rect 25780 32302 25832 32308
rect 25792 31754 25820 32302
rect 25792 31726 25912 31754
rect 25780 31680 25832 31686
rect 25780 31622 25832 31628
rect 25792 30258 25820 31622
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 25792 30054 25820 30194
rect 25780 30048 25832 30054
rect 25780 29990 25832 29996
rect 25780 29504 25832 29510
rect 25780 29446 25832 29452
rect 25608 25486 25728 25514
rect 25412 24880 25464 24886
rect 25412 24822 25464 24828
rect 25412 24744 25464 24750
rect 25412 24686 25464 24692
rect 25424 24410 25452 24686
rect 25504 24608 25556 24614
rect 25504 24550 25556 24556
rect 25516 24410 25544 24550
rect 25412 24404 25464 24410
rect 25412 24346 25464 24352
rect 25504 24404 25556 24410
rect 25504 24346 25556 24352
rect 25320 24200 25372 24206
rect 25320 24142 25372 24148
rect 25332 23798 25360 24142
rect 25320 23792 25372 23798
rect 25320 23734 25372 23740
rect 25318 23216 25374 23225
rect 25318 23151 25374 23160
rect 25332 22098 25360 23151
rect 25608 22778 25636 25486
rect 25688 22976 25740 22982
rect 25688 22918 25740 22924
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25320 22092 25372 22098
rect 25320 22034 25372 22040
rect 25700 22030 25728 22918
rect 25792 22642 25820 29446
rect 25884 28778 25912 31726
rect 25976 30734 26004 32370
rect 26056 31816 26108 31822
rect 26160 31804 26188 32982
rect 26108 31776 26188 31804
rect 26056 31758 26108 31764
rect 25964 30728 26016 30734
rect 25964 30670 26016 30676
rect 25964 30252 26016 30258
rect 26068 30240 26096 31758
rect 26148 31680 26200 31686
rect 26148 31622 26200 31628
rect 26160 30734 26188 31622
rect 26148 30728 26200 30734
rect 26148 30670 26200 30676
rect 26252 30569 26280 36518
rect 26424 36100 26476 36106
rect 26424 36042 26476 36048
rect 26332 35080 26384 35086
rect 26332 35022 26384 35028
rect 26344 32774 26372 35022
rect 26436 34610 26464 36042
rect 26516 35692 26568 35698
rect 26516 35634 26568 35640
rect 26528 35290 26556 35634
rect 26608 35488 26660 35494
rect 26608 35430 26660 35436
rect 26516 35284 26568 35290
rect 26516 35226 26568 35232
rect 26424 34604 26476 34610
rect 26424 34546 26476 34552
rect 26424 34468 26476 34474
rect 26424 34410 26476 34416
rect 26436 33930 26464 34410
rect 26424 33924 26476 33930
rect 26424 33866 26476 33872
rect 26332 32768 26384 32774
rect 26332 32710 26384 32716
rect 26528 31362 26556 35226
rect 26620 35154 26648 35430
rect 26608 35148 26660 35154
rect 26608 35090 26660 35096
rect 26700 35080 26752 35086
rect 26700 35022 26752 35028
rect 26712 34746 26740 35022
rect 26792 35012 26844 35018
rect 26792 34954 26844 34960
rect 26700 34740 26752 34746
rect 26700 34682 26752 34688
rect 26804 33561 26832 34954
rect 26976 33992 27028 33998
rect 26976 33934 27028 33940
rect 26790 33552 26846 33561
rect 26608 33516 26660 33522
rect 26790 33487 26846 33496
rect 26608 33458 26660 33464
rect 26620 33114 26648 33458
rect 26608 33108 26660 33114
rect 26608 33050 26660 33056
rect 26608 32768 26660 32774
rect 26608 32710 26660 32716
rect 26620 32065 26648 32710
rect 26700 32292 26752 32298
rect 26700 32234 26752 32240
rect 26606 32056 26662 32065
rect 26606 31991 26662 32000
rect 26606 31920 26662 31929
rect 26712 31906 26740 32234
rect 26662 31878 26740 31906
rect 26606 31855 26662 31864
rect 26712 31822 26740 31878
rect 26700 31816 26752 31822
rect 26700 31758 26752 31764
rect 26424 31340 26476 31346
rect 26528 31334 26648 31362
rect 26424 31282 26476 31288
rect 26436 31142 26464 31282
rect 26516 31272 26568 31278
rect 26516 31214 26568 31220
rect 26424 31136 26476 31142
rect 26344 31096 26424 31124
rect 26238 30560 26294 30569
rect 26238 30495 26294 30504
rect 26148 30252 26200 30258
rect 26068 30212 26148 30240
rect 25964 30194 26016 30200
rect 26148 30194 26200 30200
rect 26240 30252 26292 30258
rect 26240 30194 26292 30200
rect 25976 29753 26004 30194
rect 26056 30116 26108 30122
rect 26056 30058 26108 30064
rect 26068 29782 26096 30058
rect 26056 29776 26108 29782
rect 25962 29744 26018 29753
rect 26056 29718 26108 29724
rect 25962 29679 26018 29688
rect 26056 29640 26108 29646
rect 26056 29582 26108 29588
rect 25964 29164 26016 29170
rect 25964 29106 26016 29112
rect 25976 28994 26004 29106
rect 26068 28994 26096 29582
rect 25976 28966 26096 28994
rect 25964 28960 26016 28966
rect 25964 28902 26016 28908
rect 25884 28750 26004 28778
rect 25872 28484 25924 28490
rect 25872 28426 25924 28432
rect 25884 26874 25912 28426
rect 25976 26994 26004 28750
rect 26160 28626 26188 30194
rect 26148 28620 26200 28626
rect 26148 28562 26200 28568
rect 26252 28257 26280 30194
rect 26344 29646 26372 31096
rect 26424 31078 26476 31084
rect 26424 30728 26476 30734
rect 26424 30670 26476 30676
rect 26436 29646 26464 30670
rect 26528 30258 26556 31214
rect 26620 30734 26648 31334
rect 26804 31278 26832 33487
rect 26884 32972 26936 32978
rect 26884 32914 26936 32920
rect 26896 31754 26924 32914
rect 26988 31958 27016 33934
rect 26976 31952 27028 31958
rect 26976 31894 27028 31900
rect 26896 31726 27016 31754
rect 26792 31272 26844 31278
rect 26792 31214 26844 31220
rect 26700 31204 26752 31210
rect 26700 31146 26752 31152
rect 26608 30728 26660 30734
rect 26608 30670 26660 30676
rect 26712 30433 26740 31146
rect 26804 30802 26832 31214
rect 26792 30796 26844 30802
rect 26792 30738 26844 30744
rect 26698 30424 26754 30433
rect 26698 30359 26754 30368
rect 26608 30320 26660 30326
rect 26608 30262 26660 30268
rect 26516 30252 26568 30258
rect 26516 30194 26568 30200
rect 26620 30122 26648 30262
rect 26608 30116 26660 30122
rect 26608 30058 26660 30064
rect 26700 30048 26752 30054
rect 26700 29990 26752 29996
rect 26712 29782 26740 29990
rect 26700 29776 26752 29782
rect 26700 29718 26752 29724
rect 26332 29640 26384 29646
rect 26332 29582 26384 29588
rect 26424 29640 26476 29646
rect 26792 29640 26844 29646
rect 26424 29582 26476 29588
rect 26712 29600 26792 29628
rect 26436 29306 26464 29582
rect 26516 29504 26568 29510
rect 26516 29446 26568 29452
rect 26528 29306 26556 29446
rect 26424 29300 26476 29306
rect 26424 29242 26476 29248
rect 26516 29300 26568 29306
rect 26516 29242 26568 29248
rect 26712 29034 26740 29600
rect 26792 29582 26844 29588
rect 26884 29164 26936 29170
rect 26884 29106 26936 29112
rect 26700 29028 26752 29034
rect 26700 28970 26752 28976
rect 26238 28248 26294 28257
rect 26238 28183 26294 28192
rect 26516 27872 26568 27878
rect 26516 27814 26568 27820
rect 26056 27396 26108 27402
rect 26056 27338 26108 27344
rect 26068 27130 26096 27338
rect 26424 27328 26476 27334
rect 26424 27270 26476 27276
rect 26056 27124 26108 27130
rect 26056 27066 26108 27072
rect 26330 27024 26386 27033
rect 25964 26988 26016 26994
rect 26436 26994 26464 27270
rect 26330 26959 26386 26968
rect 26424 26988 26476 26994
rect 25964 26930 26016 26936
rect 25884 26846 26004 26874
rect 25872 26784 25924 26790
rect 25872 26726 25924 26732
rect 25884 26353 25912 26726
rect 25870 26344 25926 26353
rect 25870 26279 25926 26288
rect 25884 24818 25912 26279
rect 25976 25770 26004 26846
rect 26056 26852 26108 26858
rect 26056 26794 26108 26800
rect 26068 26382 26096 26794
rect 26148 26512 26200 26518
rect 26148 26454 26200 26460
rect 26056 26376 26108 26382
rect 26056 26318 26108 26324
rect 26056 26240 26108 26246
rect 26056 26182 26108 26188
rect 26068 26042 26096 26182
rect 26056 26036 26108 26042
rect 26056 25978 26108 25984
rect 26056 25832 26108 25838
rect 26056 25774 26108 25780
rect 25964 25764 26016 25770
rect 25964 25706 26016 25712
rect 26068 25294 26096 25774
rect 26160 25362 26188 26454
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 26252 25430 26280 26318
rect 26344 25906 26372 26959
rect 26424 26930 26476 26936
rect 26528 26926 26556 27814
rect 26712 27674 26740 28970
rect 26792 28212 26844 28218
rect 26792 28154 26844 28160
rect 26700 27668 26752 27674
rect 26700 27610 26752 27616
rect 26516 26920 26568 26926
rect 26516 26862 26568 26868
rect 26422 26480 26478 26489
rect 26422 26415 26478 26424
rect 26332 25900 26384 25906
rect 26332 25842 26384 25848
rect 26332 25764 26384 25770
rect 26332 25706 26384 25712
rect 26344 25673 26372 25706
rect 26330 25664 26386 25673
rect 26330 25599 26386 25608
rect 26436 25430 26464 26415
rect 26240 25424 26292 25430
rect 26240 25366 26292 25372
rect 26424 25424 26476 25430
rect 26424 25366 26476 25372
rect 26148 25356 26200 25362
rect 26148 25298 26200 25304
rect 26056 25288 26108 25294
rect 26056 25230 26108 25236
rect 26424 24880 26476 24886
rect 26424 24822 26476 24828
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25976 24274 26004 24550
rect 25964 24268 26016 24274
rect 25964 24210 26016 24216
rect 26436 23866 26464 24822
rect 26528 24070 26556 26862
rect 26712 26450 26740 27610
rect 26700 26444 26752 26450
rect 26700 26386 26752 26392
rect 26608 25696 26660 25702
rect 26608 25638 26660 25644
rect 26516 24064 26568 24070
rect 26516 24006 26568 24012
rect 26424 23860 26476 23866
rect 26424 23802 26476 23808
rect 25870 23760 25926 23769
rect 25870 23695 25926 23704
rect 26056 23724 26108 23730
rect 25884 23662 25912 23695
rect 26056 23666 26108 23672
rect 25872 23656 25924 23662
rect 25872 23598 25924 23604
rect 25884 23050 25912 23598
rect 26068 23322 26096 23666
rect 26056 23316 26108 23322
rect 26056 23258 26108 23264
rect 26332 23316 26384 23322
rect 26332 23258 26384 23264
rect 26056 23112 26108 23118
rect 25962 23080 26018 23089
rect 25872 23044 25924 23050
rect 26056 23054 26108 23060
rect 25962 23015 25964 23024
rect 25872 22986 25924 22992
rect 26016 23015 26018 23024
rect 25964 22986 26016 22992
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 25792 22030 25820 22578
rect 25872 22568 25924 22574
rect 25872 22510 25924 22516
rect 25884 22234 25912 22510
rect 26068 22506 26096 23054
rect 26240 22976 26292 22982
rect 26240 22918 26292 22924
rect 26252 22778 26280 22918
rect 26240 22772 26292 22778
rect 26240 22714 26292 22720
rect 26148 22636 26200 22642
rect 26148 22578 26200 22584
rect 26056 22500 26108 22506
rect 26056 22442 26108 22448
rect 25964 22432 26016 22438
rect 25964 22374 26016 22380
rect 25872 22228 25924 22234
rect 25872 22170 25924 22176
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 25780 22024 25832 22030
rect 25780 21966 25832 21972
rect 25320 21616 25372 21622
rect 25320 21558 25372 21564
rect 25332 21146 25360 21558
rect 25504 21548 25556 21554
rect 25504 21490 25556 21496
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 25516 21078 25544 21490
rect 25700 21162 25728 21966
rect 25870 21720 25926 21729
rect 25870 21655 25926 21664
rect 25884 21622 25912 21655
rect 25872 21616 25924 21622
rect 25872 21558 25924 21564
rect 25700 21134 25912 21162
rect 25504 21072 25556 21078
rect 25504 21014 25556 21020
rect 25688 21072 25740 21078
rect 25688 21014 25740 21020
rect 25318 20632 25374 20641
rect 25318 20567 25374 20576
rect 25504 20596 25556 20602
rect 25228 20460 25280 20466
rect 25228 20402 25280 20408
rect 25332 20398 25360 20567
rect 25504 20538 25556 20544
rect 25320 20392 25372 20398
rect 25320 20334 25372 20340
rect 25412 20392 25464 20398
rect 25412 20334 25464 20340
rect 25516 20346 25544 20538
rect 25332 19938 25360 20334
rect 25148 19910 25360 19938
rect 25148 19854 25176 19910
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 25228 19780 25280 19786
rect 25228 19722 25280 19728
rect 25320 19780 25372 19786
rect 25320 19722 25372 19728
rect 25240 19292 25268 19722
rect 25332 19417 25360 19722
rect 25318 19408 25374 19417
rect 25318 19343 25374 19352
rect 25424 19292 25452 20334
rect 25516 20318 25636 20346
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25516 19854 25544 20198
rect 25504 19848 25556 19854
rect 25504 19790 25556 19796
rect 25240 19264 25452 19292
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 25136 18284 25188 18290
rect 25240 18272 25268 19264
rect 25188 18244 25268 18272
rect 25412 18284 25464 18290
rect 25136 18226 25188 18232
rect 25516 18272 25544 19790
rect 25608 18630 25636 20318
rect 25700 19242 25728 21014
rect 25884 20466 25912 21134
rect 25872 20460 25924 20466
rect 25872 20402 25924 20408
rect 25872 19848 25924 19854
rect 25872 19790 25924 19796
rect 25778 19544 25834 19553
rect 25884 19514 25912 19790
rect 25778 19479 25834 19488
rect 25872 19508 25924 19514
rect 25688 19236 25740 19242
rect 25688 19178 25740 19184
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25464 18244 25544 18272
rect 25412 18226 25464 18232
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24674 17096 24730 17105
rect 24674 17031 24730 17040
rect 24584 16992 24636 16998
rect 24584 16934 24636 16940
rect 24490 16552 24546 16561
rect 24490 16487 24546 16496
rect 24504 16153 24532 16487
rect 24490 16144 24546 16153
rect 24490 16079 24546 16088
rect 24504 15706 24532 16079
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24504 15502 24532 15642
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 24124 14884 24176 14890
rect 24124 14826 24176 14832
rect 24596 14822 24624 16934
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24688 15502 24716 16050
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24688 15366 24716 15438
rect 24676 15360 24728 15366
rect 24676 15302 24728 15308
rect 24584 14816 24636 14822
rect 24584 14758 24636 14764
rect 24124 14408 24176 14414
rect 24124 14350 24176 14356
rect 24136 13938 24164 14350
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24136 13326 24164 13874
rect 24400 13796 24452 13802
rect 24400 13738 24452 13744
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24124 13320 24176 13326
rect 24124 13262 24176 13268
rect 24228 12850 24256 13670
rect 24216 12844 24268 12850
rect 24216 12786 24268 12792
rect 24124 12776 24176 12782
rect 24124 12718 24176 12724
rect 24136 11762 24164 12718
rect 24228 11762 24256 12786
rect 24308 12776 24360 12782
rect 24308 12718 24360 12724
rect 24320 12442 24348 12718
rect 24308 12436 24360 12442
rect 24308 12378 24360 12384
rect 24412 12238 24440 13738
rect 24492 13252 24544 13258
rect 24492 13194 24544 13200
rect 24504 12866 24532 13194
rect 24504 12838 24624 12866
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 24504 11778 24532 12718
rect 24412 11762 24532 11778
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24400 11756 24532 11762
rect 24452 11750 24532 11756
rect 24596 11778 24624 12838
rect 24688 12288 24716 15302
rect 24780 14890 24808 17614
rect 25148 17066 25176 18226
rect 25136 17060 25188 17066
rect 25136 17002 25188 17008
rect 25424 16726 25452 18226
rect 25700 18154 25728 19178
rect 25792 18222 25820 19479
rect 25872 19450 25924 19456
rect 25884 18902 25912 19450
rect 25872 18896 25924 18902
rect 25872 18838 25924 18844
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25688 18148 25740 18154
rect 25688 18090 25740 18096
rect 25412 16720 25464 16726
rect 25412 16662 25464 16668
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24872 16114 24900 16594
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25148 16182 25176 16390
rect 25240 16250 25268 16526
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25136 16176 25188 16182
rect 25136 16118 25188 16124
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 24952 15904 25004 15910
rect 24952 15846 25004 15852
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 24768 14884 24820 14890
rect 24768 14826 24820 14832
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 24780 12986 24808 13874
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24872 12714 24900 13262
rect 24860 12708 24912 12714
rect 24860 12650 24912 12656
rect 24768 12300 24820 12306
rect 24688 12260 24768 12288
rect 24768 12242 24820 12248
rect 24596 11762 24716 11778
rect 24780 11762 24808 12242
rect 24596 11756 24728 11762
rect 24596 11750 24676 11756
rect 24400 11698 24452 11704
rect 24676 11698 24728 11704
rect 24768 11756 24820 11762
rect 24768 11698 24820 11704
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 24136 10198 24164 11698
rect 24228 11218 24256 11698
rect 24216 11212 24268 11218
rect 24216 11154 24268 11160
rect 24412 10810 24440 11698
rect 24400 10804 24452 10810
rect 24400 10746 24452 10752
rect 24400 10600 24452 10606
rect 24400 10542 24452 10548
rect 24124 10192 24176 10198
rect 24124 10134 24176 10140
rect 24122 9888 24178 9897
rect 24122 9823 24178 9832
rect 24136 9722 24164 9823
rect 24412 9738 24440 10542
rect 24490 9888 24546 9897
rect 24546 9846 24624 9874
rect 24490 9823 24546 9832
rect 24124 9716 24176 9722
rect 24412 9710 24532 9738
rect 24124 9658 24176 9664
rect 24308 9444 24360 9450
rect 24308 9386 24360 9392
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 23938 9208 23994 9217
rect 23938 9143 23994 9152
rect 24136 8566 24164 9318
rect 24320 8634 24348 9386
rect 24400 9104 24452 9110
rect 24400 9046 24452 9052
rect 24412 8974 24440 9046
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 24308 8628 24360 8634
rect 24308 8570 24360 8576
rect 24124 8560 24176 8566
rect 24124 8502 24176 8508
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 22940 8350 23152 8378
rect 23296 8424 23348 8430
rect 23296 8366 23348 8372
rect 22940 7478 22968 8350
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23032 7954 23060 8230
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 23112 7812 23164 7818
rect 23112 7754 23164 7760
rect 23124 7546 23152 7754
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 22928 7472 22980 7478
rect 22928 7414 22980 7420
rect 22940 6390 22968 7414
rect 23308 6458 23336 8366
rect 23584 8090 23612 8434
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23584 7410 23612 8026
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 24044 7410 24072 7958
rect 24504 7410 24532 9710
rect 24596 9110 24624 9846
rect 24688 9194 24716 11698
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24780 9353 24808 11154
rect 24964 9926 24992 15846
rect 25056 13938 25084 15846
rect 25148 15473 25176 16118
rect 25240 15502 25268 16186
rect 25516 15502 25544 16458
rect 25228 15496 25280 15502
rect 25134 15464 25190 15473
rect 25228 15438 25280 15444
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25134 15399 25190 15408
rect 25516 15366 25544 15438
rect 25504 15360 25556 15366
rect 25504 15302 25556 15308
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25700 15026 25728 15302
rect 25688 15020 25740 15026
rect 25688 14962 25740 14968
rect 25596 14816 25648 14822
rect 25596 14758 25648 14764
rect 25504 14408 25556 14414
rect 25504 14350 25556 14356
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 25148 13938 25176 14214
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 25136 13932 25188 13938
rect 25136 13874 25188 13880
rect 25516 13802 25544 14350
rect 25504 13796 25556 13802
rect 25504 13738 25556 13744
rect 25608 13326 25636 14758
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25792 14006 25820 14214
rect 25780 14000 25832 14006
rect 25780 13942 25832 13948
rect 25780 13728 25832 13734
rect 25780 13670 25832 13676
rect 25792 13394 25820 13670
rect 25780 13388 25832 13394
rect 25780 13330 25832 13336
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25504 13252 25556 13258
rect 25504 13194 25556 13200
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 25148 12442 25176 12582
rect 25240 12442 25268 12718
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 25228 12436 25280 12442
rect 25228 12378 25280 12384
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 25056 11354 25084 11698
rect 25044 11348 25096 11354
rect 25044 11290 25096 11296
rect 25516 10248 25544 13194
rect 25608 12850 25636 13262
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25792 12714 25820 13126
rect 25884 12986 25912 13262
rect 25872 12980 25924 12986
rect 25872 12922 25924 12928
rect 25780 12708 25832 12714
rect 25780 12650 25832 12656
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25792 11558 25820 12038
rect 25780 11552 25832 11558
rect 25780 11494 25832 11500
rect 25792 11014 25820 11494
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25688 10260 25740 10266
rect 25516 10220 25688 10248
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24872 9722 24900 9862
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24964 9654 24992 9862
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 24766 9344 24822 9353
rect 24822 9302 24992 9330
rect 24766 9279 24822 9288
rect 24688 9166 24900 9194
rect 24872 9110 24900 9166
rect 24584 9104 24636 9110
rect 24584 9046 24636 9052
rect 24860 9104 24912 9110
rect 24860 9046 24912 9052
rect 24964 8974 24992 9302
rect 25516 9217 25544 9454
rect 25502 9208 25558 9217
rect 25502 9143 25558 9152
rect 24952 8968 25004 8974
rect 24952 8910 25004 8916
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 24584 8900 24636 8906
rect 24584 8842 24636 8848
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 24596 7410 24624 8842
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 23572 7268 23624 7274
rect 23572 7210 23624 7216
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 22928 6384 22980 6390
rect 22928 6326 22980 6332
rect 22836 5908 22888 5914
rect 22836 5850 22888 5856
rect 22940 5710 22968 6326
rect 23584 6322 23612 7210
rect 24044 6322 24072 7346
rect 24492 7200 24544 7206
rect 24492 7142 24544 7148
rect 24504 6390 24532 7142
rect 24492 6384 24544 6390
rect 24492 6326 24544 6332
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22928 5704 22980 5710
rect 22928 5646 22980 5652
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 22848 5370 22876 5510
rect 22836 5364 22888 5370
rect 22836 5306 22888 5312
rect 23032 5234 23060 6054
rect 23124 5710 23152 6258
rect 24400 6180 24452 6186
rect 24400 6122 24452 6128
rect 23204 5908 23256 5914
rect 23204 5850 23256 5856
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 23124 5234 23152 5646
rect 23216 5234 23244 5850
rect 24412 5710 24440 6122
rect 24688 5846 24716 8434
rect 25044 7812 25096 7818
rect 25044 7754 25096 7760
rect 25056 7478 25084 7754
rect 25044 7472 25096 7478
rect 25044 7414 25096 7420
rect 25148 7206 25176 8774
rect 25332 8566 25360 8842
rect 25320 8560 25372 8566
rect 25320 8502 25372 8508
rect 25424 8430 25452 8910
rect 25412 8424 25464 8430
rect 25464 8384 25544 8412
rect 25412 8366 25464 8372
rect 25320 8288 25372 8294
rect 25320 8230 25372 8236
rect 25332 7478 25360 8230
rect 25320 7472 25372 7478
rect 25320 7414 25372 7420
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 24860 7200 24912 7206
rect 24860 7142 24912 7148
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 24872 6866 24900 7142
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24964 6458 24992 6734
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 24676 5840 24728 5846
rect 25056 5794 25084 7142
rect 25240 6458 25268 7346
rect 25412 7336 25464 7342
rect 25412 7278 25464 7284
rect 25424 7002 25452 7278
rect 25412 6996 25464 7002
rect 25412 6938 25464 6944
rect 25412 6724 25464 6730
rect 25412 6666 25464 6672
rect 25320 6656 25372 6662
rect 25320 6598 25372 6604
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 25332 6390 25360 6598
rect 25320 6384 25372 6390
rect 25320 6326 25372 6332
rect 24676 5782 24728 5788
rect 24964 5778 25084 5794
rect 24952 5772 25084 5778
rect 25004 5766 25084 5772
rect 24952 5714 25004 5720
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23664 5704 23716 5710
rect 23664 5646 23716 5652
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 23584 5370 23612 5646
rect 23676 5370 23704 5646
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 23572 5364 23624 5370
rect 23572 5306 23624 5312
rect 23664 5364 23716 5370
rect 23664 5306 23716 5312
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 23112 5228 23164 5234
rect 23112 5170 23164 5176
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 21824 4616 21876 4622
rect 21822 4584 21824 4593
rect 21876 4584 21878 4593
rect 20076 4548 20128 4554
rect 20076 4490 20128 4496
rect 20536 4548 20588 4554
rect 22756 4554 22784 5170
rect 24412 5166 24440 5510
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24400 5160 24452 5166
rect 24400 5102 24452 5108
rect 23296 5092 23348 5098
rect 23296 5034 23348 5040
rect 23308 4672 23336 5034
rect 23388 5024 23440 5030
rect 23388 4966 23440 4972
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 23400 4826 23428 4966
rect 24412 4826 24440 4966
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 23480 4684 23532 4690
rect 23308 4644 23480 4672
rect 23308 4554 23336 4644
rect 23480 4626 23532 4632
rect 24688 4554 24716 5170
rect 24872 4622 24900 5306
rect 25424 5234 25452 6666
rect 25412 5228 25464 5234
rect 25412 5170 25464 5176
rect 25516 4826 25544 8384
rect 25608 6798 25636 10220
rect 25688 10202 25740 10208
rect 25792 8906 25820 10950
rect 25872 8968 25924 8974
rect 25872 8910 25924 8916
rect 25780 8900 25832 8906
rect 25780 8842 25832 8848
rect 25884 7818 25912 8910
rect 25872 7812 25924 7818
rect 25872 7754 25924 7760
rect 25596 6792 25648 6798
rect 25596 6734 25648 6740
rect 25608 6662 25636 6734
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 25504 4820 25556 4826
rect 25504 4762 25556 4768
rect 25412 4684 25464 4690
rect 25412 4626 25464 4632
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 25134 4584 25190 4593
rect 21822 4519 21878 4528
rect 22744 4548 22796 4554
rect 20536 4490 20588 4496
rect 22744 4490 22796 4496
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 24492 4548 24544 4554
rect 24676 4548 24728 4554
rect 24544 4508 24676 4536
rect 24492 4490 24544 4496
rect 25134 4519 25190 4528
rect 24676 4490 24728 4496
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 25148 4146 25176 4519
rect 25136 4140 25188 4146
rect 25228 4140 25280 4146
rect 25188 4100 25228 4128
rect 25136 4082 25188 4088
rect 25228 4082 25280 4088
rect 25424 4010 25452 4626
rect 25516 4282 25544 4762
rect 25596 4616 25648 4622
rect 25594 4584 25596 4593
rect 25648 4584 25650 4593
rect 25594 4519 25650 4528
rect 25504 4276 25556 4282
rect 25504 4218 25556 4224
rect 25412 4004 25464 4010
rect 25412 3946 25464 3952
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 25976 3058 26004 22374
rect 26068 22098 26096 22442
rect 26056 22092 26108 22098
rect 26056 22034 26108 22040
rect 26056 21548 26108 21554
rect 26056 21490 26108 21496
rect 26068 21321 26096 21490
rect 26054 21312 26110 21321
rect 26054 21247 26110 21256
rect 26056 20460 26108 20466
rect 26056 20402 26108 20408
rect 26068 20097 26096 20402
rect 26160 20330 26188 22578
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 26252 20466 26280 21966
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 26148 20324 26200 20330
rect 26148 20266 26200 20272
rect 26054 20088 26110 20097
rect 26344 20058 26372 23258
rect 26436 20058 26464 23802
rect 26620 22642 26648 25638
rect 26712 25158 26740 26386
rect 26804 25294 26832 28154
rect 26896 25498 26924 29106
rect 26884 25492 26936 25498
rect 26884 25434 26936 25440
rect 26792 25288 26844 25294
rect 26792 25230 26844 25236
rect 26700 25152 26752 25158
rect 26700 25094 26752 25100
rect 26988 24342 27016 31726
rect 27080 29034 27108 37742
rect 28000 37369 28028 37742
rect 27986 37360 28042 37369
rect 27896 37324 27948 37330
rect 27986 37295 28042 37304
rect 27896 37266 27948 37272
rect 27344 37256 27396 37262
rect 27344 37198 27396 37204
rect 27356 36174 27384 37198
rect 27620 37120 27672 37126
rect 27620 37062 27672 37068
rect 27436 36576 27488 36582
rect 27436 36518 27488 36524
rect 27252 36168 27304 36174
rect 27252 36110 27304 36116
rect 27344 36168 27396 36174
rect 27344 36110 27396 36116
rect 27264 34406 27292 36110
rect 27356 35698 27384 36110
rect 27344 35692 27396 35698
rect 27344 35634 27396 35640
rect 27448 35630 27476 36518
rect 27436 35624 27488 35630
rect 27436 35566 27488 35572
rect 27632 35086 27660 37062
rect 27804 36916 27856 36922
rect 27804 36858 27856 36864
rect 27712 36780 27764 36786
rect 27712 36722 27764 36728
rect 27344 35080 27396 35086
rect 27344 35022 27396 35028
rect 27620 35080 27672 35086
rect 27620 35022 27672 35028
rect 27252 34400 27304 34406
rect 27252 34342 27304 34348
rect 27160 33856 27212 33862
rect 27160 33798 27212 33804
rect 27172 33658 27200 33798
rect 27356 33658 27384 35022
rect 27160 33652 27212 33658
rect 27160 33594 27212 33600
rect 27344 33652 27396 33658
rect 27344 33594 27396 33600
rect 27528 32904 27580 32910
rect 27528 32846 27580 32852
rect 27252 32768 27304 32774
rect 27252 32710 27304 32716
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 27172 30938 27200 31282
rect 27160 30932 27212 30938
rect 27160 30874 27212 30880
rect 27068 29028 27120 29034
rect 27068 28970 27120 28976
rect 26976 24336 27028 24342
rect 26976 24278 27028 24284
rect 27080 23730 27108 28970
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 27172 25158 27200 25842
rect 27160 25152 27212 25158
rect 27160 25094 27212 25100
rect 27172 24857 27200 25094
rect 27158 24848 27214 24857
rect 27158 24783 27214 24792
rect 27160 23792 27212 23798
rect 27160 23734 27212 23740
rect 27068 23724 27120 23730
rect 27068 23666 27120 23672
rect 27172 23594 27200 23734
rect 27160 23588 27212 23594
rect 27160 23530 27212 23536
rect 27172 22642 27200 23530
rect 26516 22636 26568 22642
rect 26516 22578 26568 22584
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 26528 22030 26556 22578
rect 26620 22098 26648 22578
rect 26608 22092 26660 22098
rect 27264 22094 27292 32710
rect 27540 32570 27568 32846
rect 27632 32774 27660 35022
rect 27620 32768 27672 32774
rect 27620 32710 27672 32716
rect 27528 32564 27580 32570
rect 27528 32506 27580 32512
rect 27724 32502 27752 36722
rect 27816 35834 27844 36858
rect 27908 36718 27936 37266
rect 27988 37188 28040 37194
rect 27988 37130 28040 37136
rect 27896 36712 27948 36718
rect 27896 36654 27948 36660
rect 27804 35828 27856 35834
rect 27804 35770 27856 35776
rect 27816 34950 27844 35770
rect 27908 35170 27936 36654
rect 28000 36242 28028 37130
rect 28264 36780 28316 36786
rect 28264 36722 28316 36728
rect 28172 36712 28224 36718
rect 28172 36654 28224 36660
rect 27988 36236 28040 36242
rect 27988 36178 28040 36184
rect 28184 36020 28212 36654
rect 28276 36378 28304 36722
rect 28448 36576 28500 36582
rect 28448 36518 28500 36524
rect 28264 36372 28316 36378
rect 28264 36314 28316 36320
rect 28264 36168 28316 36174
rect 28316 36116 28396 36122
rect 28264 36110 28396 36116
rect 28276 36094 28396 36110
rect 28184 35992 28304 36020
rect 28276 35630 28304 35992
rect 28172 35624 28224 35630
rect 28172 35566 28224 35572
rect 28264 35624 28316 35630
rect 28264 35566 28316 35572
rect 28184 35290 28212 35566
rect 28368 35290 28396 36094
rect 28460 36009 28488 36518
rect 28552 36174 28580 38150
rect 29000 37868 29052 37874
rect 29000 37810 29052 37816
rect 28632 37324 28684 37330
rect 28632 37266 28684 37272
rect 28644 36582 28672 37266
rect 29012 36922 29040 37810
rect 29288 37262 29316 38218
rect 29472 38010 29500 38218
rect 29460 38004 29512 38010
rect 29460 37946 29512 37952
rect 29460 37800 29512 37806
rect 29460 37742 29512 37748
rect 29276 37256 29328 37262
rect 29276 37198 29328 37204
rect 29000 36916 29052 36922
rect 29000 36858 29052 36864
rect 29368 36780 29420 36786
rect 29368 36722 29420 36728
rect 29276 36644 29328 36650
rect 29276 36586 29328 36592
rect 28632 36576 28684 36582
rect 28632 36518 28684 36524
rect 28540 36168 28592 36174
rect 28540 36110 28592 36116
rect 28446 36000 28502 36009
rect 28446 35935 28502 35944
rect 28448 35624 28500 35630
rect 28448 35566 28500 35572
rect 28172 35284 28224 35290
rect 28172 35226 28224 35232
rect 28356 35284 28408 35290
rect 28356 35226 28408 35232
rect 28080 35216 28132 35222
rect 27908 35142 28028 35170
rect 28080 35158 28132 35164
rect 27896 35080 27948 35086
rect 27896 35022 27948 35028
rect 27804 34944 27856 34950
rect 27804 34886 27856 34892
rect 27804 33448 27856 33454
rect 27804 33390 27856 33396
rect 27816 32978 27844 33390
rect 27804 32972 27856 32978
rect 27804 32914 27856 32920
rect 27712 32496 27764 32502
rect 27712 32438 27764 32444
rect 27724 31754 27752 32438
rect 27908 31822 27936 35022
rect 28000 32366 28028 35142
rect 28092 35086 28120 35158
rect 28080 35080 28132 35086
rect 28080 35022 28132 35028
rect 28170 34504 28226 34513
rect 28368 34490 28396 35226
rect 28460 34649 28488 35566
rect 28552 34678 28580 36110
rect 28540 34672 28592 34678
rect 28446 34640 28502 34649
rect 28540 34614 28592 34620
rect 28446 34575 28502 34584
rect 28226 34462 28396 34490
rect 28170 34439 28226 34448
rect 28080 34400 28132 34406
rect 28080 34342 28132 34348
rect 28092 34202 28120 34342
rect 28080 34196 28132 34202
rect 28080 34138 28132 34144
rect 28448 34128 28500 34134
rect 28448 34070 28500 34076
rect 28460 33998 28488 34070
rect 28448 33992 28500 33998
rect 28448 33934 28500 33940
rect 28172 33856 28224 33862
rect 28172 33798 28224 33804
rect 28080 32836 28132 32842
rect 28080 32778 28132 32784
rect 28092 32570 28120 32778
rect 28080 32564 28132 32570
rect 28080 32506 28132 32512
rect 27988 32360 28040 32366
rect 27988 32302 28040 32308
rect 27896 31816 27948 31822
rect 27896 31758 27948 31764
rect 28184 31754 28212 33798
rect 28552 33590 28580 34614
rect 28644 33998 28672 36518
rect 29288 36378 29316 36586
rect 29276 36372 29328 36378
rect 29276 36314 29328 36320
rect 28724 36236 28776 36242
rect 28724 36178 28776 36184
rect 28736 35766 28764 36178
rect 28724 35760 28776 35766
rect 28724 35702 28776 35708
rect 28632 33992 28684 33998
rect 28632 33934 28684 33940
rect 28540 33584 28592 33590
rect 28540 33526 28592 33532
rect 28540 32972 28592 32978
rect 28540 32914 28592 32920
rect 28356 32360 28408 32366
rect 28356 32302 28408 32308
rect 28448 32360 28500 32366
rect 28448 32302 28500 32308
rect 28264 31816 28316 31822
rect 28264 31758 28316 31764
rect 27344 31748 27396 31754
rect 27344 31690 27396 31696
rect 27632 31726 27752 31754
rect 28092 31726 28212 31754
rect 27356 30190 27384 31690
rect 27632 31482 27660 31726
rect 27712 31680 27764 31686
rect 27712 31622 27764 31628
rect 27988 31680 28040 31686
rect 27988 31622 28040 31628
rect 27620 31476 27672 31482
rect 27620 31418 27672 31424
rect 27724 31278 27752 31622
rect 28000 31414 28028 31622
rect 27988 31408 28040 31414
rect 27988 31350 28040 31356
rect 27712 31272 27764 31278
rect 27712 31214 27764 31220
rect 27436 31136 27488 31142
rect 27712 31136 27764 31142
rect 27436 31078 27488 31084
rect 27710 31104 27712 31113
rect 27764 31104 27766 31113
rect 27448 30734 27476 31078
rect 27710 31039 27766 31048
rect 27620 30796 27672 30802
rect 27620 30738 27672 30744
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27344 30184 27396 30190
rect 27344 30126 27396 30132
rect 27356 29782 27384 30126
rect 27344 29776 27396 29782
rect 27344 29718 27396 29724
rect 27632 29714 27660 30738
rect 27620 29708 27672 29714
rect 27620 29650 27672 29656
rect 27344 29640 27396 29646
rect 27344 29582 27396 29588
rect 27356 29306 27384 29582
rect 27344 29300 27396 29306
rect 27344 29242 27396 29248
rect 27632 27674 27660 29650
rect 27620 27668 27672 27674
rect 27620 27610 27672 27616
rect 27436 27396 27488 27402
rect 27436 27338 27488 27344
rect 27344 26920 27396 26926
rect 27344 26862 27396 26868
rect 27356 26246 27384 26862
rect 27344 26240 27396 26246
rect 27344 26182 27396 26188
rect 27356 24886 27384 26182
rect 27344 24880 27396 24886
rect 27344 24822 27396 24828
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27356 23610 27384 24210
rect 27448 24138 27476 27338
rect 27528 25696 27580 25702
rect 27528 25638 27580 25644
rect 27540 25362 27568 25638
rect 27528 25356 27580 25362
rect 27528 25298 27580 25304
rect 27528 25220 27580 25226
rect 27528 25162 27580 25168
rect 27540 24954 27568 25162
rect 27528 24948 27580 24954
rect 27528 24890 27580 24896
rect 27540 24410 27568 24890
rect 27528 24404 27580 24410
rect 27528 24346 27580 24352
rect 27436 24132 27488 24138
rect 27436 24074 27488 24080
rect 27620 24064 27672 24070
rect 27620 24006 27672 24012
rect 27528 23724 27580 23730
rect 27528 23666 27580 23672
rect 27356 23594 27476 23610
rect 27356 23588 27488 23594
rect 27356 23582 27436 23588
rect 27356 23118 27384 23582
rect 27436 23530 27488 23536
rect 27540 23474 27568 23666
rect 27632 23594 27660 24006
rect 27724 23730 27752 31039
rect 27804 30320 27856 30326
rect 27804 30262 27856 30268
rect 27816 30122 27844 30262
rect 27804 30116 27856 30122
rect 27804 30058 27856 30064
rect 27988 30116 28040 30122
rect 27988 30058 28040 30064
rect 28000 29510 28028 30058
rect 27988 29504 28040 29510
rect 27988 29446 28040 29452
rect 27804 27328 27856 27334
rect 27804 27270 27856 27276
rect 27896 27328 27948 27334
rect 27896 27270 27948 27276
rect 27816 27130 27844 27270
rect 27804 27124 27856 27130
rect 27804 27066 27856 27072
rect 27908 26926 27936 27270
rect 27896 26920 27948 26926
rect 27896 26862 27948 26868
rect 27804 26240 27856 26246
rect 27804 26182 27856 26188
rect 27816 24750 27844 26182
rect 27894 25528 27950 25537
rect 27894 25463 27950 25472
rect 27908 25430 27936 25463
rect 27896 25424 27948 25430
rect 27896 25366 27948 25372
rect 27804 24744 27856 24750
rect 27804 24686 27856 24692
rect 27712 23724 27764 23730
rect 27712 23666 27764 23672
rect 27620 23588 27672 23594
rect 27620 23530 27672 23536
rect 27712 23588 27764 23594
rect 27712 23530 27764 23536
rect 27448 23446 27568 23474
rect 27344 23112 27396 23118
rect 27344 23054 27396 23060
rect 27448 22642 27476 23446
rect 27724 23361 27752 23530
rect 27710 23352 27766 23361
rect 27710 23287 27766 23296
rect 27528 23248 27580 23254
rect 27528 23190 27580 23196
rect 27540 22778 27568 23190
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 27724 22137 27752 22578
rect 27710 22128 27766 22137
rect 26608 22034 26660 22040
rect 26988 22066 27292 22094
rect 27528 22092 27580 22098
rect 26516 22024 26568 22030
rect 26516 21966 26568 21972
rect 26700 21684 26752 21690
rect 26700 21626 26752 21632
rect 26712 20942 26740 21626
rect 26988 21146 27016 22066
rect 27448 22052 27528 22080
rect 27448 21418 27476 22052
rect 27710 22063 27766 22072
rect 27528 22034 27580 22040
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 27620 21888 27672 21894
rect 27620 21830 27672 21836
rect 27712 21888 27764 21894
rect 27712 21830 27764 21836
rect 27804 21888 27856 21894
rect 27804 21830 27856 21836
rect 27436 21412 27488 21418
rect 27436 21354 27488 21360
rect 26976 21140 27028 21146
rect 26976 21082 27028 21088
rect 27448 21010 27476 21354
rect 27540 21146 27568 21830
rect 27528 21140 27580 21146
rect 27528 21082 27580 21088
rect 27436 21004 27488 21010
rect 27436 20946 27488 20952
rect 26700 20936 26752 20942
rect 26700 20878 26752 20884
rect 27252 20936 27304 20942
rect 27252 20878 27304 20884
rect 26712 20466 26740 20878
rect 26884 20868 26936 20874
rect 26884 20810 26936 20816
rect 26700 20460 26752 20466
rect 26700 20402 26752 20408
rect 26054 20023 26110 20032
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 26424 20052 26476 20058
rect 26424 19994 26476 20000
rect 26332 19916 26384 19922
rect 26332 19858 26384 19864
rect 26344 19825 26372 19858
rect 26712 19854 26740 20402
rect 26700 19848 26752 19854
rect 26330 19816 26386 19825
rect 26700 19790 26752 19796
rect 26330 19751 26386 19760
rect 26792 19780 26844 19786
rect 26792 19722 26844 19728
rect 26804 19174 26832 19722
rect 26792 19168 26844 19174
rect 26792 19110 26844 19116
rect 26804 18970 26832 19110
rect 26792 18964 26844 18970
rect 26792 18906 26844 18912
rect 26056 18624 26108 18630
rect 26056 18566 26108 18572
rect 26068 18290 26096 18566
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 26240 18148 26292 18154
rect 26240 18090 26292 18096
rect 26252 17814 26280 18090
rect 26516 18080 26568 18086
rect 26516 18022 26568 18028
rect 26240 17808 26292 17814
rect 26240 17750 26292 17756
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26056 16584 26108 16590
rect 26056 16526 26108 16532
rect 26068 15502 26096 16526
rect 26252 15502 26280 16594
rect 26424 16448 26476 16454
rect 26424 16390 26476 16396
rect 26436 16114 26464 16390
rect 26424 16108 26476 16114
rect 26424 16050 26476 16056
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 26068 15162 26096 15438
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 26332 15020 26384 15026
rect 26332 14962 26384 14968
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26148 14952 26200 14958
rect 26344 14929 26372 14962
rect 26148 14894 26200 14900
rect 26330 14920 26386 14929
rect 26160 13938 26188 14894
rect 26330 14855 26386 14864
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 26240 14272 26292 14278
rect 26240 14214 26292 14220
rect 26148 13932 26200 13938
rect 26148 13874 26200 13880
rect 26252 13818 26280 14214
rect 26344 14074 26372 14758
rect 26436 14618 26464 14962
rect 26424 14612 26476 14618
rect 26424 14554 26476 14560
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 26160 13790 26280 13818
rect 26160 12594 26188 13790
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26252 13394 26280 13670
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 26344 12850 26372 14010
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26160 12566 26280 12594
rect 26252 12306 26280 12566
rect 26332 12436 26384 12442
rect 26332 12378 26384 12384
rect 26344 12306 26372 12378
rect 26436 12322 26464 14554
rect 26528 13326 26556 18022
rect 26896 17882 26924 20810
rect 27264 20466 27292 20878
rect 27632 20806 27660 21830
rect 27724 21690 27752 21830
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27724 21457 27752 21490
rect 27710 21448 27766 21457
rect 27710 21383 27766 21392
rect 27710 21176 27766 21185
rect 27816 21162 27844 21830
rect 27896 21616 27948 21622
rect 27894 21584 27896 21593
rect 27948 21584 27950 21593
rect 27894 21519 27950 21528
rect 27766 21134 27844 21162
rect 27710 21111 27766 21120
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 28000 20602 28028 29446
rect 27988 20596 28040 20602
rect 27988 20538 28040 20544
rect 27252 20460 27304 20466
rect 27172 20420 27252 20448
rect 27172 19854 27200 20420
rect 27620 20460 27672 20466
rect 27252 20402 27304 20408
rect 27356 20420 27620 20448
rect 27252 20324 27304 20330
rect 27252 20266 27304 20272
rect 27264 19854 27292 20266
rect 27356 19961 27384 20420
rect 27620 20402 27672 20408
rect 27528 20324 27580 20330
rect 27528 20266 27580 20272
rect 27342 19952 27398 19961
rect 27342 19887 27398 19896
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27172 19514 27200 19790
rect 27160 19508 27212 19514
rect 27160 19450 27212 19456
rect 27068 19440 27120 19446
rect 27066 19408 27068 19417
rect 27120 19408 27122 19417
rect 27066 19343 27122 19352
rect 27172 19360 27200 19450
rect 27252 19372 27304 19378
rect 27172 19332 27252 19360
rect 27252 19314 27304 19320
rect 26884 17876 26936 17882
rect 26884 17818 26936 17824
rect 27356 17610 27384 19887
rect 27540 19446 27568 20266
rect 27618 19544 27674 19553
rect 28092 19514 28120 31726
rect 28276 30938 28304 31758
rect 28264 30932 28316 30938
rect 28264 30874 28316 30880
rect 28368 29594 28396 32302
rect 28460 30598 28488 32302
rect 28552 30682 28580 32914
rect 28644 30802 28672 33934
rect 28736 33402 28764 35702
rect 28816 34944 28868 34950
rect 28816 34886 28868 34892
rect 28828 34746 28856 34886
rect 28816 34740 28868 34746
rect 28816 34682 28868 34688
rect 28816 33856 28868 33862
rect 28816 33798 28868 33804
rect 28828 33590 28856 33798
rect 28816 33584 28868 33590
rect 28816 33526 28868 33532
rect 29184 33516 29236 33522
rect 29184 33458 29236 33464
rect 28736 33374 28856 33402
rect 28828 32910 28856 33374
rect 28816 32904 28868 32910
rect 28816 32846 28868 32852
rect 29092 32836 29144 32842
rect 29092 32778 29144 32784
rect 28724 32768 28776 32774
rect 28724 32710 28776 32716
rect 28736 32434 28764 32710
rect 28724 32428 28776 32434
rect 28724 32370 28776 32376
rect 28736 31958 28764 32370
rect 28724 31952 28776 31958
rect 28724 31894 28776 31900
rect 29104 31890 29132 32778
rect 29092 31884 29144 31890
rect 29092 31826 29144 31832
rect 29104 31754 29132 31826
rect 29012 31726 29132 31754
rect 29012 31226 29040 31726
rect 29012 31198 29132 31226
rect 29196 31210 29224 33458
rect 29276 31816 29328 31822
rect 29276 31758 29328 31764
rect 29288 31657 29316 31758
rect 29274 31648 29330 31657
rect 29274 31583 29330 31592
rect 29000 31136 29052 31142
rect 29000 31078 29052 31084
rect 28632 30796 28684 30802
rect 28632 30738 28684 30744
rect 28552 30654 28672 30682
rect 29012 30666 29040 31078
rect 28448 30592 28500 30598
rect 28500 30552 28580 30580
rect 28448 30534 28500 30540
rect 28276 29566 28396 29594
rect 28276 27878 28304 29566
rect 28356 29504 28408 29510
rect 28356 29446 28408 29452
rect 28368 29306 28396 29446
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 28264 27872 28316 27878
rect 28264 27814 28316 27820
rect 28356 27600 28408 27606
rect 28356 27542 28408 27548
rect 28172 27464 28224 27470
rect 28172 27406 28224 27412
rect 28184 26586 28212 27406
rect 28264 27328 28316 27334
rect 28264 27270 28316 27276
rect 28276 26897 28304 27270
rect 28262 26888 28318 26897
rect 28262 26823 28318 26832
rect 28264 26784 28316 26790
rect 28264 26726 28316 26732
rect 28172 26580 28224 26586
rect 28172 26522 28224 26528
rect 28276 26450 28304 26726
rect 28368 26450 28396 27542
rect 28264 26444 28316 26450
rect 28264 26386 28316 26392
rect 28356 26444 28408 26450
rect 28356 26386 28408 26392
rect 28276 25294 28304 26386
rect 28264 25288 28316 25294
rect 28264 25230 28316 25236
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28184 23798 28212 24142
rect 28172 23792 28224 23798
rect 28172 23734 28224 23740
rect 28368 22778 28396 26386
rect 28448 24200 28500 24206
rect 28448 24142 28500 24148
rect 28356 22772 28408 22778
rect 28356 22714 28408 22720
rect 28460 22234 28488 24142
rect 28264 22228 28316 22234
rect 28264 22170 28316 22176
rect 28448 22228 28500 22234
rect 28448 22170 28500 22176
rect 28276 21962 28304 22170
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 28264 21956 28316 21962
rect 28184 21916 28264 21944
rect 27618 19479 27674 19488
rect 28080 19508 28132 19514
rect 27436 19440 27488 19446
rect 27436 19382 27488 19388
rect 27528 19440 27580 19446
rect 27528 19382 27580 19388
rect 27448 18902 27476 19382
rect 27632 19378 27660 19479
rect 28080 19450 28132 19456
rect 27988 19440 28040 19446
rect 27908 19417 27988 19428
rect 27894 19408 27988 19417
rect 27620 19372 27672 19378
rect 27620 19314 27672 19320
rect 27804 19372 27856 19378
rect 27950 19400 27988 19408
rect 27988 19382 28040 19388
rect 27894 19343 27950 19352
rect 28080 19372 28132 19378
rect 27804 19314 27856 19320
rect 28080 19314 28132 19320
rect 27436 18896 27488 18902
rect 27436 18838 27488 18844
rect 27710 17776 27766 17785
rect 27710 17711 27712 17720
rect 27764 17711 27766 17720
rect 27712 17682 27764 17688
rect 27816 17678 27844 19314
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 27896 18080 27948 18086
rect 27896 18022 27948 18028
rect 27908 17678 27936 18022
rect 28000 17882 28028 18226
rect 27988 17876 28040 17882
rect 27988 17818 28040 17824
rect 28092 17762 28120 19314
rect 28184 19310 28212 21916
rect 28264 21898 28316 21904
rect 28262 19408 28318 19417
rect 28262 19343 28264 19352
rect 28316 19343 28318 19352
rect 28264 19314 28316 19320
rect 28172 19304 28224 19310
rect 28172 19246 28224 19252
rect 28184 18290 28212 19246
rect 28460 18630 28488 21966
rect 28552 21894 28580 30552
rect 28644 29170 28672 30654
rect 29000 30660 29052 30666
rect 29000 30602 29052 30608
rect 29104 30394 29132 31198
rect 29184 31204 29236 31210
rect 29184 31146 29236 31152
rect 29092 30388 29144 30394
rect 29092 30330 29144 30336
rect 28724 29776 28776 29782
rect 28724 29718 28776 29724
rect 28736 29646 28764 29718
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 28724 29640 28776 29646
rect 28724 29582 28776 29588
rect 29012 29306 29040 29650
rect 29000 29300 29052 29306
rect 29000 29242 29052 29248
rect 28632 29164 28684 29170
rect 28632 29106 28684 29112
rect 28644 27130 28672 29106
rect 29092 28756 29144 28762
rect 29092 28698 29144 28704
rect 29104 28218 29132 28698
rect 29092 28212 29144 28218
rect 29092 28154 29144 28160
rect 28816 27872 28868 27878
rect 28736 27832 28816 27860
rect 28632 27124 28684 27130
rect 28632 27066 28684 27072
rect 28632 25832 28684 25838
rect 28632 25774 28684 25780
rect 28644 25294 28672 25774
rect 28632 25288 28684 25294
rect 28632 25230 28684 25236
rect 28736 22094 28764 27832
rect 28816 27814 28868 27820
rect 29092 27532 29144 27538
rect 29092 27474 29144 27480
rect 29000 26852 29052 26858
rect 29000 26794 29052 26800
rect 29012 26382 29040 26794
rect 29000 26376 29052 26382
rect 29000 26318 29052 26324
rect 28908 25424 28960 25430
rect 28908 25366 28960 25372
rect 28816 24812 28868 24818
rect 28816 24754 28868 24760
rect 28828 23866 28856 24754
rect 28816 23860 28868 23866
rect 28816 23802 28868 23808
rect 28920 23798 28948 25366
rect 29104 25362 29132 27474
rect 29196 27470 29224 31146
rect 29288 29782 29316 31583
rect 29276 29776 29328 29782
rect 29276 29718 29328 29724
rect 29276 29504 29328 29510
rect 29276 29446 29328 29452
rect 29288 29306 29316 29446
rect 29276 29300 29328 29306
rect 29276 29242 29328 29248
rect 29276 28960 29328 28966
rect 29276 28902 29328 28908
rect 29288 28762 29316 28902
rect 29276 28756 29328 28762
rect 29276 28698 29328 28704
rect 29184 27464 29236 27470
rect 29184 27406 29236 27412
rect 29276 26512 29328 26518
rect 29276 26454 29328 26460
rect 29184 26308 29236 26314
rect 29184 26250 29236 26256
rect 29092 25356 29144 25362
rect 29092 25298 29144 25304
rect 29092 25152 29144 25158
rect 29092 25094 29144 25100
rect 29104 24954 29132 25094
rect 29092 24948 29144 24954
rect 29092 24890 29144 24896
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 28908 23792 28960 23798
rect 28908 23734 28960 23740
rect 28736 22066 28856 22094
rect 28724 22024 28776 22030
rect 28724 21966 28776 21972
rect 28540 21888 28592 21894
rect 28540 21830 28592 21836
rect 28736 21418 28764 21966
rect 28828 21622 28856 22066
rect 29012 21894 29040 24550
rect 29092 22024 29144 22030
rect 29092 21966 29144 21972
rect 29000 21888 29052 21894
rect 29000 21830 29052 21836
rect 28816 21616 28868 21622
rect 28816 21558 28868 21564
rect 28724 21412 28776 21418
rect 28724 21354 28776 21360
rect 28724 20392 28776 20398
rect 28724 20334 28776 20340
rect 28816 20392 28868 20398
rect 28816 20334 28868 20340
rect 28632 20324 28684 20330
rect 28632 20266 28684 20272
rect 28644 20058 28672 20266
rect 28632 20052 28684 20058
rect 28632 19994 28684 20000
rect 28736 19922 28764 20334
rect 28828 20058 28856 20334
rect 28908 20256 28960 20262
rect 28908 20198 28960 20204
rect 28920 20058 28948 20198
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28908 20052 28960 20058
rect 28908 19994 28960 20000
rect 28998 19952 29054 19961
rect 28724 19916 28776 19922
rect 28998 19887 29054 19896
rect 28724 19858 28776 19864
rect 28540 19780 28592 19786
rect 28540 19722 28592 19728
rect 28552 19378 28580 19722
rect 28736 19514 28764 19858
rect 29012 19836 29040 19887
rect 28966 19808 29040 19836
rect 28966 19718 28994 19808
rect 28954 19712 29006 19718
rect 29104 19689 29132 21966
rect 29196 21350 29224 26250
rect 29288 26081 29316 26454
rect 29274 26072 29330 26081
rect 29274 26007 29330 26016
rect 29380 23322 29408 36722
rect 29472 36718 29500 37742
rect 29564 37330 29592 38286
rect 29656 38010 29684 38286
rect 29644 38004 29696 38010
rect 29644 37946 29696 37952
rect 29552 37324 29604 37330
rect 29552 37266 29604 37272
rect 29460 36712 29512 36718
rect 29460 36654 29512 36660
rect 29564 35222 29592 37266
rect 29644 36712 29696 36718
rect 29644 36654 29696 36660
rect 29656 35494 29684 36654
rect 29644 35488 29696 35494
rect 29644 35430 29696 35436
rect 29552 35216 29604 35222
rect 29552 35158 29604 35164
rect 29644 34400 29696 34406
rect 29644 34342 29696 34348
rect 29656 33862 29684 34342
rect 29644 33856 29696 33862
rect 29644 33798 29696 33804
rect 29458 33144 29514 33153
rect 29458 33079 29514 33088
rect 29552 33108 29604 33114
rect 29472 24206 29500 33079
rect 29552 33050 29604 33056
rect 29564 31822 29592 33050
rect 29552 31816 29604 31822
rect 29552 31758 29604 31764
rect 29552 31680 29604 31686
rect 29552 31622 29604 31628
rect 29564 31142 29592 31622
rect 29644 31340 29696 31346
rect 29644 31282 29696 31288
rect 29552 31136 29604 31142
rect 29552 31078 29604 31084
rect 29656 30938 29684 31282
rect 29644 30932 29696 30938
rect 29644 30874 29696 30880
rect 29644 29640 29696 29646
rect 29644 29582 29696 29588
rect 29552 29504 29604 29510
rect 29552 29446 29604 29452
rect 29460 24200 29512 24206
rect 29460 24142 29512 24148
rect 29368 23316 29420 23322
rect 29368 23258 29420 23264
rect 29184 21344 29236 21350
rect 29184 21286 29236 21292
rect 29460 20936 29512 20942
rect 29460 20878 29512 20884
rect 29368 19780 29420 19786
rect 29368 19722 29420 19728
rect 29184 19712 29236 19718
rect 28954 19654 29006 19660
rect 29090 19680 29146 19689
rect 29184 19654 29236 19660
rect 29090 19615 29146 19624
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28540 19372 28592 19378
rect 28540 19314 28592 19320
rect 28448 18624 28500 18630
rect 28448 18566 28500 18572
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28632 18216 28684 18222
rect 28632 18158 28684 18164
rect 28092 17746 28304 17762
rect 28092 17740 28316 17746
rect 28092 17734 28264 17740
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 27896 17672 27948 17678
rect 27896 17614 27948 17620
rect 27988 17672 28040 17678
rect 27988 17614 28040 17620
rect 27344 17604 27396 17610
rect 27344 17546 27396 17552
rect 27816 17202 27844 17614
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 27160 15972 27212 15978
rect 27160 15914 27212 15920
rect 27344 15972 27396 15978
rect 27344 15914 27396 15920
rect 27172 15570 27200 15914
rect 27356 15706 27384 15914
rect 27436 15904 27488 15910
rect 27436 15846 27488 15852
rect 27344 15700 27396 15706
rect 27344 15642 27396 15648
rect 27448 15570 27476 15846
rect 27160 15564 27212 15570
rect 27436 15564 27488 15570
rect 27212 15524 27292 15552
rect 27160 15506 27212 15512
rect 27068 15496 27120 15502
rect 27068 15438 27120 15444
rect 27080 14278 27108 15438
rect 27160 15020 27212 15026
rect 27160 14962 27212 14968
rect 27172 14414 27200 14962
rect 27160 14408 27212 14414
rect 27160 14350 27212 14356
rect 27068 14272 27120 14278
rect 27068 14214 27120 14220
rect 27080 13938 27108 14214
rect 27264 14074 27292 15524
rect 27436 15506 27488 15512
rect 27436 15428 27488 15434
rect 27436 15370 27488 15376
rect 27344 15360 27396 15366
rect 27344 15302 27396 15308
rect 27356 15162 27384 15302
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 27252 14068 27304 14074
rect 27252 14010 27304 14016
rect 27068 13932 27120 13938
rect 27068 13874 27120 13880
rect 27252 13796 27304 13802
rect 27252 13738 27304 13744
rect 26700 13728 26752 13734
rect 26700 13670 26752 13676
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 26516 13320 26568 13326
rect 26568 13280 26648 13308
rect 26516 13262 26568 13268
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26528 12850 26556 13126
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 26620 12442 26648 13280
rect 26712 13258 26740 13670
rect 26976 13456 27028 13462
rect 26976 13398 27028 13404
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26700 13252 26752 13258
rect 26700 13194 26752 13200
rect 26712 12986 26740 13194
rect 26700 12980 26752 12986
rect 26700 12922 26752 12928
rect 26804 12442 26832 13262
rect 26884 12776 26936 12782
rect 26884 12718 26936 12724
rect 26608 12436 26660 12442
rect 26608 12378 26660 12384
rect 26792 12436 26844 12442
rect 26792 12378 26844 12384
rect 26240 12300 26292 12306
rect 26240 12242 26292 12248
rect 26332 12300 26384 12306
rect 26436 12294 26740 12322
rect 26332 12242 26384 12248
rect 26252 11150 26280 12242
rect 26344 11218 26372 12242
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26436 11694 26464 12174
rect 26608 12096 26660 12102
rect 26608 12038 26660 12044
rect 26620 11830 26648 12038
rect 26608 11824 26660 11830
rect 26608 11766 26660 11772
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 26436 11150 26464 11630
rect 26608 11280 26660 11286
rect 26608 11222 26660 11228
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26424 11144 26476 11150
rect 26424 11086 26476 11092
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26424 10124 26476 10130
rect 26424 10066 26476 10072
rect 26148 10056 26200 10062
rect 26148 9998 26200 10004
rect 26160 9586 26188 9998
rect 26332 9988 26384 9994
rect 26332 9930 26384 9936
rect 26148 9580 26200 9586
rect 26148 9522 26200 9528
rect 26344 8922 26372 9930
rect 26252 8894 26372 8922
rect 26252 8090 26280 8894
rect 26332 8832 26384 8838
rect 26330 8800 26332 8809
rect 26384 8800 26386 8809
rect 26330 8735 26386 8744
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 26252 7478 26280 8026
rect 26344 7478 26372 8735
rect 26436 7546 26464 10066
rect 26528 9382 26556 11086
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26528 9042 26556 9318
rect 26620 9178 26648 11222
rect 26608 9172 26660 9178
rect 26608 9114 26660 9120
rect 26516 9036 26568 9042
rect 26516 8978 26568 8984
rect 26516 8832 26568 8838
rect 26516 8774 26568 8780
rect 26528 8498 26556 8774
rect 26516 8492 26568 8498
rect 26516 8434 26568 8440
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 26608 7540 26660 7546
rect 26608 7482 26660 7488
rect 26240 7472 26292 7478
rect 26240 7414 26292 7420
rect 26332 7472 26384 7478
rect 26332 7414 26384 7420
rect 26620 7002 26648 7482
rect 26712 7206 26740 12294
rect 26896 11558 26924 12718
rect 26884 11552 26936 11558
rect 26884 11494 26936 11500
rect 26988 11132 27016 13398
rect 27172 13326 27200 13670
rect 27068 13320 27120 13326
rect 27068 13262 27120 13268
rect 27160 13320 27212 13326
rect 27160 13262 27212 13268
rect 27080 11286 27108 13262
rect 27160 12232 27212 12238
rect 27160 12174 27212 12180
rect 27172 11898 27200 12174
rect 27160 11892 27212 11898
rect 27160 11834 27212 11840
rect 27160 11620 27212 11626
rect 27160 11562 27212 11568
rect 27068 11280 27120 11286
rect 27068 11222 27120 11228
rect 27068 11144 27120 11150
rect 26988 11104 27068 11132
rect 27068 11086 27120 11092
rect 26792 11008 26844 11014
rect 26792 10950 26844 10956
rect 27068 11008 27120 11014
rect 27068 10950 27120 10956
rect 26804 10674 26832 10950
rect 26792 10668 26844 10674
rect 26792 10610 26844 10616
rect 27080 9586 27108 10950
rect 27172 9674 27200 11562
rect 27264 10674 27292 13738
rect 27448 11830 27476 15370
rect 27618 15192 27674 15201
rect 27896 15156 27948 15162
rect 27618 15127 27620 15136
rect 27672 15127 27674 15136
rect 27620 15098 27672 15104
rect 27816 15116 27896 15144
rect 27816 15026 27844 15116
rect 27896 15098 27948 15104
rect 27804 15020 27856 15026
rect 27804 14962 27856 14968
rect 27804 14000 27856 14006
rect 27804 13942 27856 13948
rect 27816 13530 27844 13942
rect 28000 13818 28028 17614
rect 28092 16998 28120 17734
rect 28264 17682 28316 17688
rect 28644 17678 28672 18158
rect 28908 18148 28960 18154
rect 28908 18090 28960 18096
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 28632 17672 28684 17678
rect 28632 17614 28684 17620
rect 28172 17604 28224 17610
rect 28172 17546 28224 17552
rect 28184 17066 28212 17546
rect 28368 17338 28396 17614
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28632 17264 28684 17270
rect 28632 17206 28684 17212
rect 28644 17116 28672 17206
rect 28276 17088 28672 17116
rect 28172 17060 28224 17066
rect 28172 17002 28224 17008
rect 28080 16992 28132 16998
rect 28080 16934 28132 16940
rect 28080 16448 28132 16454
rect 28080 16390 28132 16396
rect 28092 15502 28120 16390
rect 28080 15496 28132 15502
rect 28080 15438 28132 15444
rect 28092 13938 28120 15438
rect 28172 14952 28224 14958
rect 28172 14894 28224 14900
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 28000 13790 28120 13818
rect 27804 13524 27856 13530
rect 27804 13466 27856 13472
rect 27618 13424 27674 13433
rect 27618 13359 27674 13368
rect 27632 11898 27660 13359
rect 27804 12300 27856 12306
rect 27804 12242 27856 12248
rect 27620 11892 27672 11898
rect 27620 11834 27672 11840
rect 27436 11824 27488 11830
rect 27436 11766 27488 11772
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27356 11286 27384 11698
rect 27528 11620 27580 11626
rect 27528 11562 27580 11568
rect 27436 11552 27488 11558
rect 27436 11494 27488 11500
rect 27448 11286 27476 11494
rect 27344 11280 27396 11286
rect 27344 11222 27396 11228
rect 27436 11280 27488 11286
rect 27436 11222 27488 11228
rect 27540 10674 27568 11562
rect 27632 11218 27660 11834
rect 27816 11830 27844 12242
rect 27804 11824 27856 11830
rect 27804 11766 27856 11772
rect 27988 11824 28040 11830
rect 27988 11766 28040 11772
rect 27710 11656 27766 11665
rect 27710 11591 27766 11600
rect 27896 11620 27948 11626
rect 27724 11558 27752 11591
rect 27896 11562 27948 11568
rect 27712 11552 27764 11558
rect 27712 11494 27764 11500
rect 27620 11212 27672 11218
rect 27620 11154 27672 11160
rect 27724 11132 27752 11494
rect 27804 11144 27856 11150
rect 27724 11104 27804 11132
rect 27804 11086 27856 11092
rect 27620 11008 27672 11014
rect 27620 10950 27672 10956
rect 27632 10810 27660 10950
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27908 10577 27936 11562
rect 28000 11558 28028 11766
rect 27988 11552 28040 11558
rect 27988 11494 28040 11500
rect 28000 11150 28028 11494
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 27894 10568 27950 10577
rect 27894 10503 27950 10512
rect 27896 10464 27948 10470
rect 27896 10406 27948 10412
rect 27986 10432 28042 10441
rect 27908 10130 27936 10406
rect 28092 10418 28120 13790
rect 28184 13530 28212 14894
rect 28172 13524 28224 13530
rect 28172 13466 28224 13472
rect 28172 12776 28224 12782
rect 28172 12718 28224 12724
rect 28184 10810 28212 12718
rect 28172 10804 28224 10810
rect 28172 10746 28224 10752
rect 28172 10532 28224 10538
rect 28172 10474 28224 10480
rect 28042 10390 28120 10418
rect 27986 10367 28042 10376
rect 28184 10130 28212 10474
rect 27896 10124 27948 10130
rect 27896 10066 27948 10072
rect 28172 10124 28224 10130
rect 28172 10066 28224 10072
rect 27896 9988 27948 9994
rect 27896 9930 27948 9936
rect 27344 9716 27396 9722
rect 27172 9664 27344 9674
rect 27172 9658 27396 9664
rect 27172 9646 27384 9658
rect 27356 9586 27384 9646
rect 27068 9580 27120 9586
rect 27068 9522 27120 9528
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27712 9580 27764 9586
rect 27712 9522 27764 9528
rect 26792 8968 26844 8974
rect 26976 8968 27028 8974
rect 26882 8936 26938 8945
rect 26844 8916 26882 8922
rect 26792 8910 26882 8916
rect 26804 8894 26882 8910
rect 26976 8910 27028 8916
rect 26882 8871 26938 8880
rect 26988 8634 27016 8910
rect 26976 8628 27028 8634
rect 26976 8570 27028 8576
rect 27080 8430 27108 9522
rect 27252 9172 27304 9178
rect 27252 9114 27304 9120
rect 27160 9104 27212 9110
rect 27160 9046 27212 9052
rect 27172 8974 27200 9046
rect 27264 8974 27292 9114
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 27252 8968 27304 8974
rect 27252 8910 27304 8916
rect 27724 8906 27752 9522
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 27712 8900 27764 8906
rect 27712 8842 27764 8848
rect 27620 8492 27672 8498
rect 27448 8452 27620 8480
rect 26792 8424 26844 8430
rect 26792 8366 26844 8372
rect 27068 8424 27120 8430
rect 27068 8366 27120 8372
rect 26700 7200 26752 7206
rect 26700 7142 26752 7148
rect 26608 6996 26660 7002
rect 26608 6938 26660 6944
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26068 6322 26096 6734
rect 26056 6316 26108 6322
rect 26056 6258 26108 6264
rect 26068 5098 26096 6258
rect 26252 5234 26280 6734
rect 26804 6254 26832 8366
rect 27344 7812 27396 7818
rect 27344 7754 27396 7760
rect 27356 7478 27384 7754
rect 27344 7472 27396 7478
rect 27344 7414 27396 7420
rect 26976 6792 27028 6798
rect 26976 6734 27028 6740
rect 26792 6248 26844 6254
rect 26792 6190 26844 6196
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26988 5166 27016 6734
rect 27448 6662 27476 8452
rect 27620 8434 27672 8440
rect 27528 8356 27580 8362
rect 27528 8298 27580 8304
rect 27540 7546 27568 8298
rect 27724 7546 27752 8842
rect 27816 8809 27844 8978
rect 27802 8800 27858 8809
rect 27802 8735 27858 8744
rect 27804 8356 27856 8362
rect 27804 8298 27856 8304
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27712 7540 27764 7546
rect 27712 7482 27764 7488
rect 27436 6656 27488 6662
rect 27436 6598 27488 6604
rect 27632 6254 27660 7482
rect 27712 7200 27764 7206
rect 27712 7142 27764 7148
rect 27724 6798 27752 7142
rect 27816 6866 27844 8298
rect 27908 6934 27936 9930
rect 28080 9376 28132 9382
rect 28080 9318 28132 9324
rect 28092 9042 28120 9318
rect 28080 9036 28132 9042
rect 28080 8978 28132 8984
rect 27988 8968 28040 8974
rect 27986 8936 27988 8945
rect 28040 8936 28042 8945
rect 27986 8871 28042 8880
rect 28276 7342 28304 17088
rect 28356 15360 28408 15366
rect 28356 15302 28408 15308
rect 28368 14618 28396 15302
rect 28446 15192 28502 15201
rect 28446 15127 28502 15136
rect 28460 15026 28488 15127
rect 28722 15056 28778 15065
rect 28448 15020 28500 15026
rect 28778 15000 28856 15008
rect 28722 14991 28724 15000
rect 28448 14962 28500 14968
rect 28776 14980 28856 15000
rect 28724 14962 28776 14968
rect 28538 14920 28594 14929
rect 28448 14884 28500 14890
rect 28538 14855 28540 14864
rect 28448 14826 28500 14832
rect 28592 14855 28594 14864
rect 28540 14826 28592 14832
rect 28356 14612 28408 14618
rect 28356 14554 28408 14560
rect 28460 14074 28488 14826
rect 28828 14822 28856 14980
rect 28816 14816 28868 14822
rect 28816 14758 28868 14764
rect 28448 14068 28500 14074
rect 28448 14010 28500 14016
rect 28816 13932 28868 13938
rect 28816 13874 28868 13880
rect 28540 13728 28592 13734
rect 28540 13670 28592 13676
rect 28356 13456 28408 13462
rect 28356 13398 28408 13404
rect 28368 10674 28396 13398
rect 28552 13326 28580 13670
rect 28540 13320 28592 13326
rect 28540 13262 28592 13268
rect 28448 13184 28500 13190
rect 28448 13126 28500 13132
rect 28460 12102 28488 13126
rect 28828 12102 28856 13874
rect 28920 13190 28948 18090
rect 29104 16402 29132 19615
rect 29196 19514 29224 19654
rect 29184 19508 29236 19514
rect 29184 19450 29236 19456
rect 29380 19378 29408 19722
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 29472 18358 29500 20878
rect 29564 20466 29592 29446
rect 29656 27538 29684 29582
rect 29748 27878 29776 38762
rect 33060 38554 33088 38898
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35636 38554 35664 38898
rect 37646 38856 37702 38865
rect 37646 38791 37648 38800
rect 37700 38791 37702 38800
rect 37922 38856 37978 38865
rect 37922 38791 37978 38800
rect 37648 38762 37700 38768
rect 37936 38554 37964 38791
rect 33048 38548 33100 38554
rect 33048 38490 33100 38496
rect 35624 38548 35676 38554
rect 35624 38490 35676 38496
rect 37924 38548 37976 38554
rect 37924 38490 37976 38496
rect 32680 38412 32732 38418
rect 32680 38354 32732 38360
rect 31668 38344 31720 38350
rect 31668 38286 31720 38292
rect 30380 38208 30432 38214
rect 30380 38150 30432 38156
rect 30392 37942 30420 38150
rect 30380 37936 30432 37942
rect 30380 37878 30432 37884
rect 30392 37176 30420 37878
rect 31208 37868 31260 37874
rect 31208 37810 31260 37816
rect 30932 37664 30984 37670
rect 30932 37606 30984 37612
rect 30944 37330 30972 37606
rect 30932 37324 30984 37330
rect 30932 37266 30984 37272
rect 30472 37188 30524 37194
rect 30392 37148 30472 37176
rect 30472 37130 30524 37136
rect 30012 37120 30064 37126
rect 30012 37062 30064 37068
rect 30024 36922 30052 37062
rect 31220 36922 31248 37810
rect 31680 37806 31708 38286
rect 31668 37800 31720 37806
rect 31668 37742 31720 37748
rect 32588 37256 32640 37262
rect 32588 37198 32640 37204
rect 31484 37188 31536 37194
rect 31484 37130 31536 37136
rect 31496 36922 31524 37130
rect 32496 37120 32548 37126
rect 32496 37062 32548 37068
rect 32508 36922 32536 37062
rect 30012 36916 30064 36922
rect 30012 36858 30064 36864
rect 31208 36916 31260 36922
rect 31208 36858 31260 36864
rect 31484 36916 31536 36922
rect 31484 36858 31536 36864
rect 32496 36916 32548 36922
rect 32496 36858 32548 36864
rect 30024 36310 30052 36858
rect 30656 36712 30708 36718
rect 30656 36654 30708 36660
rect 32220 36712 32272 36718
rect 32220 36654 32272 36660
rect 30668 36378 30696 36654
rect 32232 36378 32260 36654
rect 30656 36372 30708 36378
rect 30656 36314 30708 36320
rect 32220 36372 32272 36378
rect 32220 36314 32272 36320
rect 30012 36304 30064 36310
rect 30012 36246 30064 36252
rect 29828 36100 29880 36106
rect 29828 36042 29880 36048
rect 29840 35698 29868 36042
rect 30024 35698 30052 36246
rect 30472 35760 30524 35766
rect 30472 35702 30524 35708
rect 29828 35692 29880 35698
rect 29828 35634 29880 35640
rect 30012 35692 30064 35698
rect 30012 35634 30064 35640
rect 29840 33998 29868 35634
rect 29920 35488 29972 35494
rect 29920 35430 29972 35436
rect 30104 35488 30156 35494
rect 30104 35430 30156 35436
rect 29932 35290 29960 35430
rect 29920 35284 29972 35290
rect 29920 35226 29972 35232
rect 29932 34134 29960 35226
rect 29920 34128 29972 34134
rect 29920 34070 29972 34076
rect 29828 33992 29880 33998
rect 29828 33934 29880 33940
rect 29840 31822 29868 33934
rect 29932 31906 29960 34070
rect 29932 31878 30052 31906
rect 30024 31822 30052 31878
rect 29828 31816 29880 31822
rect 30012 31816 30064 31822
rect 29880 31776 29960 31804
rect 29828 31758 29880 31764
rect 29828 30252 29880 30258
rect 29828 30194 29880 30200
rect 29840 29753 29868 30194
rect 29932 30054 29960 31776
rect 30012 31758 30064 31764
rect 30116 30682 30144 35430
rect 30380 35080 30432 35086
rect 30380 35022 30432 35028
rect 30288 32904 30340 32910
rect 30288 32846 30340 32852
rect 30196 32768 30248 32774
rect 30196 32710 30248 32716
rect 30208 30841 30236 32710
rect 30300 31890 30328 32846
rect 30288 31884 30340 31890
rect 30288 31826 30340 31832
rect 30392 31754 30420 35022
rect 30484 33998 30512 35702
rect 30668 34406 30696 36314
rect 30840 36100 30892 36106
rect 30840 36042 30892 36048
rect 30748 36032 30800 36038
rect 30748 35974 30800 35980
rect 30760 35834 30788 35974
rect 30748 35828 30800 35834
rect 30748 35770 30800 35776
rect 30852 35018 30880 36042
rect 32600 35766 32628 37198
rect 32588 35760 32640 35766
rect 32588 35702 32640 35708
rect 31392 35692 31444 35698
rect 31392 35634 31444 35640
rect 31024 35488 31076 35494
rect 31024 35430 31076 35436
rect 31036 35154 31064 35430
rect 31024 35148 31076 35154
rect 31024 35090 31076 35096
rect 30840 35012 30892 35018
rect 30840 34954 30892 34960
rect 30852 34474 30880 34954
rect 31404 34746 31432 35634
rect 31484 35624 31536 35630
rect 31484 35566 31536 35572
rect 30932 34740 30984 34746
rect 30932 34682 30984 34688
rect 31392 34740 31444 34746
rect 31392 34682 31444 34688
rect 30840 34468 30892 34474
rect 30840 34410 30892 34416
rect 30564 34400 30616 34406
rect 30564 34342 30616 34348
rect 30656 34400 30708 34406
rect 30944 34354 30972 34682
rect 31300 34468 31352 34474
rect 31300 34410 31352 34416
rect 30656 34342 30708 34348
rect 30576 33998 30604 34342
rect 30852 34326 30972 34354
rect 30852 34202 30880 34326
rect 30840 34196 30892 34202
rect 30840 34138 30892 34144
rect 30852 33998 30880 34138
rect 30472 33992 30524 33998
rect 30472 33934 30524 33940
rect 30564 33992 30616 33998
rect 30564 33934 30616 33940
rect 30840 33992 30892 33998
rect 30840 33934 30892 33940
rect 30484 33114 30512 33934
rect 31312 33114 31340 34410
rect 31496 33998 31524 35566
rect 32496 35012 32548 35018
rect 32496 34954 32548 34960
rect 31668 34944 31720 34950
rect 31668 34886 31720 34892
rect 31576 34604 31628 34610
rect 31576 34546 31628 34552
rect 31484 33992 31536 33998
rect 31484 33934 31536 33940
rect 30472 33108 30524 33114
rect 30472 33050 30524 33056
rect 30656 33108 30708 33114
rect 30656 33050 30708 33056
rect 31300 33108 31352 33114
rect 31300 33050 31352 33056
rect 30668 32366 30696 33050
rect 30932 32904 30984 32910
rect 30932 32846 30984 32852
rect 31208 32904 31260 32910
rect 31208 32846 31260 32852
rect 30840 32428 30892 32434
rect 30840 32370 30892 32376
rect 30656 32360 30708 32366
rect 30656 32302 30708 32308
rect 30392 31726 30512 31754
rect 30380 31680 30432 31686
rect 30380 31622 30432 31628
rect 30392 31482 30420 31622
rect 30380 31476 30432 31482
rect 30380 31418 30432 31424
rect 30194 30832 30250 30841
rect 30194 30767 30250 30776
rect 30024 30654 30144 30682
rect 29920 30048 29972 30054
rect 29920 29990 29972 29996
rect 29826 29744 29882 29753
rect 29826 29679 29882 29688
rect 29840 29646 29868 29679
rect 30024 29646 30052 30654
rect 30380 29776 30432 29782
rect 30380 29718 30432 29724
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 30196 29640 30248 29646
rect 30196 29582 30248 29588
rect 29828 29504 29880 29510
rect 29828 29446 29880 29452
rect 29736 27872 29788 27878
rect 29736 27814 29788 27820
rect 29840 27690 29868 29446
rect 30012 29096 30064 29102
rect 30012 29038 30064 29044
rect 30024 28626 30052 29038
rect 30208 28966 30236 29582
rect 30196 28960 30248 28966
rect 30248 28920 30328 28948
rect 30196 28902 30248 28908
rect 30012 28620 30064 28626
rect 30012 28562 30064 28568
rect 30104 28620 30156 28626
rect 30104 28562 30156 28568
rect 29918 27976 29974 27985
rect 29918 27911 29974 27920
rect 29748 27662 29868 27690
rect 29644 27532 29696 27538
rect 29644 27474 29696 27480
rect 29644 27328 29696 27334
rect 29644 27270 29696 27276
rect 29656 27130 29684 27270
rect 29644 27124 29696 27130
rect 29644 27066 29696 27072
rect 29748 27010 29776 27662
rect 29828 27328 29880 27334
rect 29828 27270 29880 27276
rect 29840 27130 29868 27270
rect 29828 27124 29880 27130
rect 29828 27066 29880 27072
rect 29656 26982 29776 27010
rect 29656 26042 29684 26982
rect 29736 26920 29788 26926
rect 29736 26862 29788 26868
rect 29644 26036 29696 26042
rect 29644 25978 29696 25984
rect 29748 25922 29776 26862
rect 29656 25894 29776 25922
rect 29656 24886 29684 25894
rect 29644 24880 29696 24886
rect 29644 24822 29696 24828
rect 29736 24744 29788 24750
rect 29736 24686 29788 24692
rect 29748 24206 29776 24686
rect 29932 24206 29960 27911
rect 30012 27464 30064 27470
rect 30012 27406 30064 27412
rect 30024 26586 30052 27406
rect 30012 26580 30064 26586
rect 30012 26522 30064 26528
rect 30116 26450 30144 28562
rect 30196 28416 30248 28422
rect 30196 28358 30248 28364
rect 30208 28014 30236 28358
rect 30196 28008 30248 28014
rect 30196 27950 30248 27956
rect 30104 26444 30156 26450
rect 30104 26386 30156 26392
rect 30012 26376 30064 26382
rect 30012 26318 30064 26324
rect 30024 25702 30052 26318
rect 30104 26036 30156 26042
rect 30104 25978 30156 25984
rect 30012 25696 30064 25702
rect 30012 25638 30064 25644
rect 30116 25226 30144 25978
rect 30104 25220 30156 25226
rect 30104 25162 30156 25168
rect 30116 24954 30144 25162
rect 30104 24948 30156 24954
rect 30104 24890 30156 24896
rect 30116 24342 30144 24890
rect 30208 24614 30236 27950
rect 30300 25702 30328 28920
rect 30392 28558 30420 29718
rect 30380 28552 30432 28558
rect 30380 28494 30432 28500
rect 30392 27470 30420 28494
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 30380 27328 30432 27334
rect 30380 27270 30432 27276
rect 30392 26790 30420 27270
rect 30380 26784 30432 26790
rect 30380 26726 30432 26732
rect 30484 26382 30512 31726
rect 30748 31680 30800 31686
rect 30748 31622 30800 31628
rect 30654 30832 30710 30841
rect 30654 30767 30656 30776
rect 30708 30767 30710 30776
rect 30656 30738 30708 30744
rect 30656 30320 30708 30326
rect 30656 30262 30708 30268
rect 30564 30048 30616 30054
rect 30564 29990 30616 29996
rect 30576 29646 30604 29990
rect 30564 29640 30616 29646
rect 30564 29582 30616 29588
rect 30576 29345 30604 29582
rect 30668 29578 30696 30262
rect 30760 29646 30788 31622
rect 30852 30598 30880 32370
rect 30944 32298 30972 32846
rect 31220 32570 31248 32846
rect 31208 32564 31260 32570
rect 31208 32506 31260 32512
rect 30932 32292 30984 32298
rect 30932 32234 30984 32240
rect 31496 31822 31524 33934
rect 31588 33590 31616 34546
rect 31680 34542 31708 34886
rect 31668 34536 31720 34542
rect 31668 34478 31720 34484
rect 31680 33862 31708 34478
rect 31668 33856 31720 33862
rect 31668 33798 31720 33804
rect 32220 33856 32272 33862
rect 32220 33798 32272 33804
rect 31576 33584 31628 33590
rect 31576 33526 31628 33532
rect 32128 32768 32180 32774
rect 32128 32710 32180 32716
rect 32140 32434 32168 32710
rect 32232 32434 32260 33798
rect 32508 32910 32536 34954
rect 32496 32904 32548 32910
rect 32496 32846 32548 32852
rect 32600 32502 32628 35702
rect 32588 32496 32640 32502
rect 32588 32438 32640 32444
rect 32128 32428 32180 32434
rect 32128 32370 32180 32376
rect 32220 32428 32272 32434
rect 32220 32370 32272 32376
rect 32140 32026 32168 32370
rect 32312 32360 32364 32366
rect 32312 32302 32364 32308
rect 32128 32020 32180 32026
rect 32128 31962 32180 31968
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 31024 30796 31076 30802
rect 31024 30738 31076 30744
rect 30930 30696 30986 30705
rect 30930 30631 30932 30640
rect 30984 30631 30986 30640
rect 30932 30602 30984 30608
rect 30840 30592 30892 30598
rect 30840 30534 30892 30540
rect 31036 30326 31064 30738
rect 31300 30592 31352 30598
rect 31300 30534 31352 30540
rect 31024 30320 31076 30326
rect 31024 30262 31076 30268
rect 31312 30258 31340 30534
rect 31300 30252 31352 30258
rect 31300 30194 31352 30200
rect 30840 30184 30892 30190
rect 30840 30126 30892 30132
rect 30748 29640 30800 29646
rect 30748 29582 30800 29588
rect 30656 29572 30708 29578
rect 30656 29514 30708 29520
rect 30562 29336 30618 29345
rect 30562 29271 30618 29280
rect 30576 28472 30604 29271
rect 30852 29238 30880 30126
rect 31312 29646 31340 30194
rect 31024 29640 31076 29646
rect 31024 29582 31076 29588
rect 31300 29640 31352 29646
rect 31300 29582 31352 29588
rect 30932 29504 30984 29510
rect 30932 29446 30984 29452
rect 30944 29306 30972 29446
rect 30932 29300 30984 29306
rect 30932 29242 30984 29248
rect 30840 29232 30892 29238
rect 31036 29186 31064 29582
rect 31116 29572 31168 29578
rect 31116 29514 31168 29520
rect 30840 29174 30892 29180
rect 30944 29158 31064 29186
rect 30656 28484 30708 28490
rect 30576 28444 30656 28472
rect 30656 28426 30708 28432
rect 30668 27470 30696 28426
rect 30944 28422 30972 29158
rect 31128 29034 31156 29514
rect 31496 29170 31524 31758
rect 32036 31680 32088 31686
rect 32036 31622 32088 31628
rect 31668 31340 31720 31346
rect 31668 31282 31720 31288
rect 31680 30802 31708 31282
rect 31944 31272 31996 31278
rect 31944 31214 31996 31220
rect 31668 30796 31720 30802
rect 31668 30738 31720 30744
rect 31956 30734 31984 31214
rect 31944 30728 31996 30734
rect 31944 30670 31996 30676
rect 32048 30258 32076 31622
rect 32324 30258 32352 32302
rect 32692 31754 32720 38354
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 37832 37120 37884 37126
rect 37832 37062 37884 37068
rect 37844 36825 37872 37062
rect 37830 36816 37886 36825
rect 33692 36780 33744 36786
rect 37830 36751 37886 36760
rect 33692 36722 33744 36728
rect 33140 36576 33192 36582
rect 33140 36518 33192 36524
rect 33152 36038 33180 36518
rect 33140 36032 33192 36038
rect 33140 35974 33192 35980
rect 32772 35488 32824 35494
rect 32772 35430 32824 35436
rect 32784 35290 32812 35430
rect 32772 35284 32824 35290
rect 32772 35226 32824 35232
rect 32772 34536 32824 34542
rect 32772 34478 32824 34484
rect 32600 31726 32720 31754
rect 32496 30728 32548 30734
rect 32496 30670 32548 30676
rect 32508 30258 32536 30670
rect 32036 30252 32088 30258
rect 32036 30194 32088 30200
rect 32312 30252 32364 30258
rect 32312 30194 32364 30200
rect 32496 30252 32548 30258
rect 32496 30194 32548 30200
rect 31668 29640 31720 29646
rect 31574 29608 31630 29617
rect 31668 29582 31720 29588
rect 31574 29543 31630 29552
rect 31588 29306 31616 29543
rect 31680 29306 31708 29582
rect 31576 29300 31628 29306
rect 31576 29242 31628 29248
rect 31668 29300 31720 29306
rect 31668 29242 31720 29248
rect 32324 29170 32352 30194
rect 31484 29164 31536 29170
rect 31484 29106 31536 29112
rect 32312 29164 32364 29170
rect 32312 29106 32364 29112
rect 31116 29028 31168 29034
rect 31116 28970 31168 28976
rect 31496 28558 31524 29106
rect 32404 28960 32456 28966
rect 32404 28902 32456 28908
rect 31576 28688 31628 28694
rect 31576 28630 31628 28636
rect 31484 28552 31536 28558
rect 31484 28494 31536 28500
rect 30932 28416 30984 28422
rect 30932 28358 30984 28364
rect 31116 28416 31168 28422
rect 31116 28358 31168 28364
rect 31484 28416 31536 28422
rect 31588 28404 31616 28630
rect 32416 28626 32444 28902
rect 32404 28620 32456 28626
rect 32404 28562 32456 28568
rect 31760 28552 31812 28558
rect 31760 28494 31812 28500
rect 31536 28376 31616 28404
rect 31484 28358 31536 28364
rect 30944 27470 30972 28358
rect 30656 27464 30708 27470
rect 30656 27406 30708 27412
rect 30932 27464 30984 27470
rect 30932 27406 30984 27412
rect 30472 26376 30524 26382
rect 30470 26344 30472 26353
rect 30524 26344 30526 26353
rect 30470 26279 30526 26288
rect 30668 25838 30696 27406
rect 30944 26450 30972 27406
rect 30932 26444 30984 26450
rect 30932 26386 30984 26392
rect 30656 25832 30708 25838
rect 30656 25774 30708 25780
rect 30288 25696 30340 25702
rect 30288 25638 30340 25644
rect 30300 25158 30328 25638
rect 30932 25288 30984 25294
rect 30932 25230 30984 25236
rect 30288 25152 30340 25158
rect 30288 25094 30340 25100
rect 30300 24682 30328 25094
rect 30944 24886 30972 25230
rect 30932 24880 30984 24886
rect 30932 24822 30984 24828
rect 31128 24818 31156 28358
rect 31496 28218 31524 28358
rect 31772 28218 31800 28494
rect 31944 28484 31996 28490
rect 31944 28426 31996 28432
rect 31956 28218 31984 28426
rect 31484 28212 31536 28218
rect 31484 28154 31536 28160
rect 31760 28212 31812 28218
rect 31760 28154 31812 28160
rect 31944 28212 31996 28218
rect 31944 28154 31996 28160
rect 31760 27328 31812 27334
rect 31760 27270 31812 27276
rect 31576 27124 31628 27130
rect 31576 27066 31628 27072
rect 31392 26784 31444 26790
rect 31392 26726 31444 26732
rect 31404 26450 31432 26726
rect 31392 26444 31444 26450
rect 31392 26386 31444 26392
rect 31588 26314 31616 27066
rect 31668 26988 31720 26994
rect 31668 26930 31720 26936
rect 31300 26308 31352 26314
rect 31300 26250 31352 26256
rect 31576 26308 31628 26314
rect 31576 26250 31628 26256
rect 31312 26042 31340 26250
rect 31574 26072 31630 26081
rect 31300 26036 31352 26042
rect 31680 26042 31708 26930
rect 31574 26007 31576 26016
rect 31300 25978 31352 25984
rect 31628 26007 31630 26016
rect 31668 26036 31720 26042
rect 31576 25978 31628 25984
rect 31668 25978 31720 25984
rect 31392 25968 31444 25974
rect 31390 25936 31392 25945
rect 31444 25936 31446 25945
rect 31772 25906 31800 27270
rect 32496 26444 32548 26450
rect 32496 26386 32548 26392
rect 32508 26081 32536 26386
rect 32494 26072 32550 26081
rect 32494 26007 32496 26016
rect 32548 26007 32550 26016
rect 32496 25978 32548 25984
rect 31390 25871 31446 25880
rect 31760 25900 31812 25906
rect 31760 25842 31812 25848
rect 31852 25492 31904 25498
rect 31852 25434 31904 25440
rect 31300 25152 31352 25158
rect 31300 25094 31352 25100
rect 31116 24812 31168 24818
rect 31116 24754 31168 24760
rect 30288 24676 30340 24682
rect 30288 24618 30340 24624
rect 30196 24608 30248 24614
rect 30196 24550 30248 24556
rect 31208 24608 31260 24614
rect 31208 24550 31260 24556
rect 31220 24410 31248 24550
rect 31208 24404 31260 24410
rect 31208 24346 31260 24352
rect 30104 24336 30156 24342
rect 30104 24278 30156 24284
rect 29736 24200 29788 24206
rect 29736 24142 29788 24148
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 30196 24064 30248 24070
rect 30196 24006 30248 24012
rect 29736 23112 29788 23118
rect 29736 23054 29788 23060
rect 29920 23112 29972 23118
rect 29920 23054 29972 23060
rect 29748 22438 29776 23054
rect 29932 22778 29960 23054
rect 30012 23044 30064 23050
rect 30012 22986 30064 22992
rect 29920 22772 29972 22778
rect 29920 22714 29972 22720
rect 29736 22432 29788 22438
rect 29736 22374 29788 22380
rect 29748 21622 29776 22374
rect 30024 22098 30052 22986
rect 30208 22642 30236 24006
rect 30196 22636 30248 22642
rect 30196 22578 30248 22584
rect 30656 22432 30708 22438
rect 30656 22374 30708 22380
rect 30012 22092 30064 22098
rect 30012 22034 30064 22040
rect 30024 21842 30052 22034
rect 30564 22024 30616 22030
rect 30564 21966 30616 21972
rect 29932 21814 30052 21842
rect 30380 21888 30432 21894
rect 30380 21830 30432 21836
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 29932 21690 29960 21814
rect 30392 21690 30420 21830
rect 29920 21684 29972 21690
rect 29920 21626 29972 21632
rect 30380 21684 30432 21690
rect 30380 21626 30432 21632
rect 29736 21616 29788 21622
rect 29736 21558 29788 21564
rect 29644 21344 29696 21350
rect 29644 21286 29696 21292
rect 29552 20460 29604 20466
rect 29552 20402 29604 20408
rect 29564 19922 29592 20402
rect 29656 20398 29684 21286
rect 30484 20942 30512 21830
rect 30576 21554 30604 21966
rect 30564 21548 30616 21554
rect 30564 21490 30616 21496
rect 30668 21010 30696 22374
rect 31024 22160 31076 22166
rect 30852 22108 31024 22114
rect 30852 22102 31076 22108
rect 30852 22086 31064 22102
rect 30656 21004 30708 21010
rect 30656 20946 30708 20952
rect 30380 20936 30432 20942
rect 30380 20878 30432 20884
rect 30472 20936 30524 20942
rect 30472 20878 30524 20884
rect 30196 20800 30248 20806
rect 30196 20742 30248 20748
rect 29644 20392 29696 20398
rect 29644 20334 29696 20340
rect 29552 19916 29604 19922
rect 29552 19858 29604 19864
rect 29656 19854 29684 20334
rect 29736 20052 29788 20058
rect 29736 19994 29788 20000
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29552 19712 29604 19718
rect 29552 19654 29604 19660
rect 29564 19514 29592 19654
rect 29748 19514 29776 19994
rect 29828 19848 29880 19854
rect 29828 19790 29880 19796
rect 29840 19514 29868 19790
rect 30208 19786 30236 20742
rect 30392 20466 30420 20878
rect 30668 20466 30696 20946
rect 30380 20460 30432 20466
rect 30380 20402 30432 20408
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30196 19780 30248 19786
rect 30196 19722 30248 19728
rect 30392 19514 30420 20402
rect 30656 20324 30708 20330
rect 30656 20266 30708 20272
rect 30668 20058 30696 20266
rect 30656 20052 30708 20058
rect 30656 19994 30708 20000
rect 30654 19952 30710 19961
rect 30748 19916 30800 19922
rect 30710 19896 30748 19904
rect 30654 19887 30748 19896
rect 30668 19876 30748 19887
rect 30748 19858 30800 19864
rect 29552 19508 29604 19514
rect 29552 19450 29604 19456
rect 29736 19508 29788 19514
rect 29736 19450 29788 19456
rect 29828 19508 29880 19514
rect 29828 19450 29880 19456
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 29552 19372 29604 19378
rect 29552 19314 29604 19320
rect 29460 18352 29512 18358
rect 29460 18294 29512 18300
rect 29564 18086 29592 19314
rect 29644 19168 29696 19174
rect 29644 19110 29696 19116
rect 29552 18080 29604 18086
rect 29552 18022 29604 18028
rect 29184 17536 29236 17542
rect 29184 17478 29236 17484
rect 29196 17338 29224 17478
rect 29184 17332 29236 17338
rect 29184 17274 29236 17280
rect 29656 17202 29684 19110
rect 30748 18624 30800 18630
rect 30748 18566 30800 18572
rect 30380 18352 30432 18358
rect 30378 18320 30380 18329
rect 30432 18320 30434 18329
rect 30378 18255 30434 18264
rect 29920 18216 29972 18222
rect 29840 18176 29920 18204
rect 29840 17814 29868 18176
rect 29920 18158 29972 18164
rect 30760 18170 30788 18566
rect 30852 18290 30880 22086
rect 31116 21956 31168 21962
rect 31116 21898 31168 21904
rect 31128 21554 31156 21898
rect 31116 21548 31168 21554
rect 31116 21490 31168 21496
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30944 21146 30972 21286
rect 30932 21140 30984 21146
rect 30932 21082 30984 21088
rect 30944 20466 30972 21082
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 31116 20460 31168 20466
rect 31116 20402 31168 20408
rect 31128 19417 31156 20402
rect 31208 20256 31260 20262
rect 31208 20198 31260 20204
rect 31220 19922 31248 20198
rect 31208 19916 31260 19922
rect 31208 19858 31260 19864
rect 31114 19408 31170 19417
rect 31114 19343 31170 19352
rect 31024 18624 31076 18630
rect 31024 18566 31076 18572
rect 31036 18290 31064 18566
rect 30840 18284 30892 18290
rect 30840 18226 30892 18232
rect 31024 18284 31076 18290
rect 31024 18226 31076 18232
rect 30760 18142 30880 18170
rect 29920 18080 29972 18086
rect 29920 18022 29972 18028
rect 29828 17808 29880 17814
rect 29828 17750 29880 17756
rect 29736 17672 29788 17678
rect 29736 17614 29788 17620
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29196 16794 29224 17138
rect 29276 16992 29328 16998
rect 29276 16934 29328 16940
rect 29368 16992 29420 16998
rect 29368 16934 29420 16940
rect 29184 16788 29236 16794
rect 29184 16730 29236 16736
rect 29288 16522 29316 16934
rect 29380 16726 29408 16934
rect 29368 16720 29420 16726
rect 29368 16662 29420 16668
rect 29276 16516 29328 16522
rect 29276 16458 29328 16464
rect 29104 16374 29316 16402
rect 29184 16244 29236 16250
rect 29184 16186 29236 16192
rect 29196 16153 29224 16186
rect 29182 16144 29238 16153
rect 29092 16108 29144 16114
rect 29182 16079 29238 16088
rect 29092 16050 29144 16056
rect 29104 15502 29132 16050
rect 29092 15496 29144 15502
rect 29092 15438 29144 15444
rect 29184 14544 29236 14550
rect 29184 14486 29236 14492
rect 29196 14074 29224 14486
rect 29288 14278 29316 16374
rect 29644 16176 29696 16182
rect 29642 16144 29644 16153
rect 29696 16144 29698 16153
rect 29642 16079 29698 16088
rect 29460 16040 29512 16046
rect 29460 15982 29512 15988
rect 29368 15904 29420 15910
rect 29368 15846 29420 15852
rect 29276 14272 29328 14278
rect 29276 14214 29328 14220
rect 29184 14068 29236 14074
rect 29184 14010 29236 14016
rect 29196 13938 29224 14010
rect 29184 13932 29236 13938
rect 29184 13874 29236 13880
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 29012 13530 29040 13806
rect 29276 13796 29328 13802
rect 29276 13738 29328 13744
rect 29000 13524 29052 13530
rect 29000 13466 29052 13472
rect 29184 13524 29236 13530
rect 29184 13466 29236 13472
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 29000 12708 29052 12714
rect 29000 12650 29052 12656
rect 29092 12708 29144 12714
rect 29092 12650 29144 12656
rect 28448 12096 28500 12102
rect 28448 12038 28500 12044
rect 28816 12096 28868 12102
rect 28816 12038 28868 12044
rect 28460 10742 28488 12038
rect 28828 11762 28856 12038
rect 29012 11762 29040 12650
rect 29104 11898 29132 12650
rect 29092 11892 29144 11898
rect 29092 11834 29144 11840
rect 28816 11756 28868 11762
rect 28816 11698 28868 11704
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29196 11354 29224 13466
rect 29288 13326 29316 13738
rect 29276 13320 29328 13326
rect 29276 13262 29328 13268
rect 29380 11898 29408 15846
rect 29472 15706 29500 15982
rect 29460 15700 29512 15706
rect 29460 15642 29512 15648
rect 29460 13728 29512 13734
rect 29460 13670 29512 13676
rect 29472 13326 29500 13670
rect 29460 13320 29512 13326
rect 29460 13262 29512 13268
rect 29644 13184 29696 13190
rect 29644 13126 29696 13132
rect 29656 12986 29684 13126
rect 29644 12980 29696 12986
rect 29644 12922 29696 12928
rect 29748 12442 29776 17614
rect 29932 14958 29960 18022
rect 30288 17808 30340 17814
rect 30024 17756 30288 17762
rect 30024 17750 30340 17756
rect 30024 17734 30328 17750
rect 29920 14952 29972 14958
rect 29920 14894 29972 14900
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 29368 11892 29420 11898
rect 29368 11834 29420 11840
rect 29736 11756 29788 11762
rect 29736 11698 29788 11704
rect 29184 11348 29236 11354
rect 29184 11290 29236 11296
rect 29644 11144 29696 11150
rect 29644 11086 29696 11092
rect 28448 10736 28500 10742
rect 28448 10678 28500 10684
rect 29092 10736 29144 10742
rect 29092 10678 29144 10684
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 28816 10668 28868 10674
rect 28816 10610 28868 10616
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 28368 10062 28396 10610
rect 28630 10432 28686 10441
rect 28630 10367 28686 10376
rect 28448 10260 28500 10266
rect 28448 10202 28500 10208
rect 28356 10056 28408 10062
rect 28356 9998 28408 10004
rect 28460 8974 28488 10202
rect 28448 8968 28500 8974
rect 28448 8910 28500 8916
rect 28540 7404 28592 7410
rect 28540 7346 28592 7352
rect 28264 7336 28316 7342
rect 28264 7278 28316 7284
rect 28080 7268 28132 7274
rect 28080 7210 28132 7216
rect 27896 6928 27948 6934
rect 27896 6870 27948 6876
rect 27804 6860 27856 6866
rect 27804 6802 27856 6808
rect 27712 6792 27764 6798
rect 27712 6734 27764 6740
rect 27988 6792 28040 6798
rect 27988 6734 28040 6740
rect 28000 6458 28028 6734
rect 28092 6730 28120 7210
rect 28552 6866 28580 7346
rect 28448 6860 28500 6866
rect 28448 6802 28500 6808
rect 28540 6860 28592 6866
rect 28540 6802 28592 6808
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 28264 6792 28316 6798
rect 28264 6734 28316 6740
rect 28080 6724 28132 6730
rect 28080 6666 28132 6672
rect 27988 6452 28040 6458
rect 27988 6394 28040 6400
rect 27804 6316 27856 6322
rect 27804 6258 27856 6264
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 27436 6180 27488 6186
rect 27436 6122 27488 6128
rect 27448 5914 27476 6122
rect 27632 6118 27660 6190
rect 27816 6118 27844 6258
rect 27620 6112 27672 6118
rect 27620 6054 27672 6060
rect 27804 6112 27856 6118
rect 27804 6054 27856 6060
rect 27436 5908 27488 5914
rect 27436 5850 27488 5856
rect 27632 5370 27660 6054
rect 27620 5364 27672 5370
rect 27620 5306 27672 5312
rect 27620 5228 27672 5234
rect 27620 5170 27672 5176
rect 27712 5228 27764 5234
rect 27712 5170 27764 5176
rect 26976 5160 27028 5166
rect 26976 5102 27028 5108
rect 26056 5092 26108 5098
rect 26056 5034 26108 5040
rect 26068 4826 26096 5034
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 26988 4690 27016 5102
rect 27632 4826 27660 5170
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 26976 4684 27028 4690
rect 26976 4626 27028 4632
rect 26332 4616 26384 4622
rect 26332 4558 26384 4564
rect 26344 4078 26372 4558
rect 27724 4486 27752 5170
rect 27896 4752 27948 4758
rect 27896 4694 27948 4700
rect 27712 4480 27764 4486
rect 27712 4422 27764 4428
rect 27908 4146 27936 4694
rect 28092 4690 28120 6666
rect 28184 6458 28212 6734
rect 28172 6452 28224 6458
rect 28172 6394 28224 6400
rect 28276 5166 28304 6734
rect 28356 6656 28408 6662
rect 28356 6598 28408 6604
rect 28368 5846 28396 6598
rect 28356 5840 28408 5846
rect 28356 5782 28408 5788
rect 28460 5302 28488 6802
rect 28644 6780 28672 10367
rect 28724 10056 28776 10062
rect 28724 9998 28776 10004
rect 28736 9586 28764 9998
rect 28724 9580 28776 9586
rect 28724 9522 28776 9528
rect 28828 9330 28856 10610
rect 28908 10192 28960 10198
rect 29012 10146 29040 10610
rect 29104 10198 29132 10678
rect 28960 10140 29040 10146
rect 28908 10134 29040 10140
rect 29092 10192 29144 10198
rect 29092 10134 29144 10140
rect 28920 10118 29040 10134
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 28920 9926 28948 9998
rect 29012 9994 29040 10118
rect 29000 9988 29052 9994
rect 29000 9930 29052 9936
rect 28908 9920 28960 9926
rect 28908 9862 28960 9868
rect 28920 9586 28948 9862
rect 28908 9580 28960 9586
rect 28908 9522 28960 9528
rect 28736 9302 28856 9330
rect 28736 7002 28764 9302
rect 29104 8838 29132 10134
rect 29656 9586 29684 11086
rect 29748 9586 29776 11698
rect 29828 11688 29880 11694
rect 29828 11630 29880 11636
rect 29644 9580 29696 9586
rect 29644 9522 29696 9528
rect 29736 9580 29788 9586
rect 29736 9522 29788 9528
rect 29736 9376 29788 9382
rect 29736 9318 29788 9324
rect 29748 9178 29776 9318
rect 29736 9172 29788 9178
rect 29736 9114 29788 9120
rect 29840 9110 29868 11630
rect 29184 9104 29236 9110
rect 29184 9046 29236 9052
rect 29828 9104 29880 9110
rect 29828 9046 29880 9052
rect 28816 8832 28868 8838
rect 28816 8774 28868 8780
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 29000 8832 29052 8838
rect 29000 8774 29052 8780
rect 29092 8832 29144 8838
rect 29092 8774 29144 8780
rect 28724 6996 28776 7002
rect 28724 6938 28776 6944
rect 28828 6798 28856 8774
rect 28920 8634 28948 8774
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 29012 8566 29040 8774
rect 29000 8560 29052 8566
rect 29000 8502 29052 8508
rect 29012 8294 29040 8502
rect 29000 8288 29052 8294
rect 29000 8230 29052 8236
rect 29000 7948 29052 7954
rect 29000 7890 29052 7896
rect 29012 7410 29040 7890
rect 29196 7410 29224 9046
rect 29368 8968 29420 8974
rect 29368 8910 29420 8916
rect 29276 8900 29328 8906
rect 29276 8842 29328 8848
rect 29288 8090 29316 8842
rect 29380 8430 29408 8910
rect 29368 8424 29420 8430
rect 29368 8366 29420 8372
rect 29644 8288 29696 8294
rect 29644 8230 29696 8236
rect 29276 8084 29328 8090
rect 29276 8026 29328 8032
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 29184 7404 29236 7410
rect 29184 7346 29236 7352
rect 28908 6996 28960 7002
rect 28908 6938 28960 6944
rect 28724 6792 28776 6798
rect 28644 6752 28724 6780
rect 28724 6734 28776 6740
rect 28816 6792 28868 6798
rect 28816 6734 28868 6740
rect 28920 6118 28948 6938
rect 28908 6112 28960 6118
rect 28908 6054 28960 6060
rect 29196 5778 29224 7346
rect 29288 5846 29316 8026
rect 29656 7546 29684 8230
rect 29932 7954 29960 14894
rect 30024 12850 30052 17734
rect 30104 17672 30156 17678
rect 30104 17614 30156 17620
rect 30288 17672 30340 17678
rect 30288 17614 30340 17620
rect 30116 17134 30144 17614
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30208 17338 30236 17478
rect 30196 17332 30248 17338
rect 30196 17274 30248 17280
rect 30104 17128 30156 17134
rect 30104 17070 30156 17076
rect 30300 16998 30328 17614
rect 30288 16992 30340 16998
rect 30288 16934 30340 16940
rect 30196 16584 30248 16590
rect 30196 16526 30248 16532
rect 30288 16584 30340 16590
rect 30288 16526 30340 16532
rect 30656 16584 30708 16590
rect 30656 16526 30708 16532
rect 30208 16250 30236 16526
rect 30196 16244 30248 16250
rect 30196 16186 30248 16192
rect 30300 16182 30328 16526
rect 30668 16454 30696 16526
rect 30656 16448 30708 16454
rect 30656 16390 30708 16396
rect 30748 16448 30800 16454
rect 30748 16390 30800 16396
rect 30760 16250 30788 16390
rect 30748 16244 30800 16250
rect 30748 16186 30800 16192
rect 30288 16176 30340 16182
rect 30288 16118 30340 16124
rect 30104 15904 30156 15910
rect 30380 15904 30432 15910
rect 30104 15846 30156 15852
rect 30208 15852 30380 15858
rect 30208 15846 30432 15852
rect 30116 13870 30144 15846
rect 30208 15830 30420 15846
rect 30208 14385 30236 15830
rect 30760 15706 30788 16186
rect 30852 16130 30880 18142
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 30944 16250 30972 16526
rect 30932 16244 30984 16250
rect 30932 16186 30984 16192
rect 30852 16102 30972 16130
rect 30748 15700 30800 15706
rect 30748 15642 30800 15648
rect 30288 15428 30340 15434
rect 30288 15370 30340 15376
rect 30300 14906 30328 15370
rect 30656 15360 30708 15366
rect 30656 15302 30708 15308
rect 30668 15026 30696 15302
rect 30656 15020 30708 15026
rect 30656 14962 30708 14968
rect 30840 15020 30892 15026
rect 30840 14962 30892 14968
rect 30564 14952 30616 14958
rect 30300 14890 30512 14906
rect 30564 14894 30616 14900
rect 30300 14884 30524 14890
rect 30300 14878 30472 14884
rect 30472 14826 30524 14832
rect 30576 14770 30604 14894
rect 30392 14742 30604 14770
rect 30194 14376 30250 14385
rect 30194 14311 30250 14320
rect 30392 14278 30420 14742
rect 30668 14482 30696 14962
rect 30748 14884 30800 14890
rect 30748 14826 30800 14832
rect 30656 14476 30708 14482
rect 30656 14418 30708 14424
rect 30196 14272 30248 14278
rect 30196 14214 30248 14220
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30104 13864 30156 13870
rect 30104 13806 30156 13812
rect 30012 12844 30064 12850
rect 30012 12786 30064 12792
rect 30012 12640 30064 12646
rect 30012 12582 30064 12588
rect 30024 12238 30052 12582
rect 30012 12232 30064 12238
rect 30012 12174 30064 12180
rect 30208 11642 30236 14214
rect 30392 13938 30420 14214
rect 30380 13932 30432 13938
rect 30380 13874 30432 13880
rect 30472 13864 30524 13870
rect 30472 13806 30524 13812
rect 30288 13456 30340 13462
rect 30288 13398 30340 13404
rect 30300 12782 30328 13398
rect 30380 12844 30432 12850
rect 30380 12786 30432 12792
rect 30288 12776 30340 12782
rect 30288 12718 30340 12724
rect 30392 12102 30420 12786
rect 30484 12238 30512 13806
rect 30668 12850 30696 14418
rect 30760 14346 30788 14826
rect 30852 14482 30880 14962
rect 30840 14476 30892 14482
rect 30840 14418 30892 14424
rect 30748 14340 30800 14346
rect 30748 14282 30800 14288
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 30852 13938 30880 14010
rect 30840 13932 30892 13938
rect 30840 13874 30892 13880
rect 30748 13796 30800 13802
rect 30748 13738 30800 13744
rect 30656 12844 30708 12850
rect 30656 12786 30708 12792
rect 30472 12232 30524 12238
rect 30524 12192 30604 12220
rect 30472 12174 30524 12180
rect 30380 12096 30432 12102
rect 30380 12038 30432 12044
rect 30472 12096 30524 12102
rect 30472 12038 30524 12044
rect 30392 11898 30420 12038
rect 30380 11892 30432 11898
rect 30380 11834 30432 11840
rect 30484 11762 30512 12038
rect 30288 11756 30340 11762
rect 30288 11698 30340 11704
rect 30472 11756 30524 11762
rect 30472 11698 30524 11704
rect 30024 11614 30236 11642
rect 30024 9489 30052 11614
rect 30300 11558 30328 11698
rect 30288 11552 30340 11558
rect 30288 11494 30340 11500
rect 30380 11552 30432 11558
rect 30380 11494 30432 11500
rect 30392 11354 30420 11494
rect 30104 11348 30156 11354
rect 30104 11290 30156 11296
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 30116 9586 30144 11290
rect 30484 11218 30512 11698
rect 30472 11212 30524 11218
rect 30472 11154 30524 11160
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30208 11014 30236 11086
rect 30196 11008 30248 11014
rect 30196 10950 30248 10956
rect 30300 10674 30328 11086
rect 30288 10668 30340 10674
rect 30288 10610 30340 10616
rect 30194 10160 30250 10169
rect 30194 10095 30250 10104
rect 30208 10062 30236 10095
rect 30196 10056 30248 10062
rect 30196 9998 30248 10004
rect 30104 9580 30156 9586
rect 30104 9522 30156 9528
rect 30010 9480 30066 9489
rect 30010 9415 30066 9424
rect 30116 8974 30144 9522
rect 30196 9512 30248 9518
rect 30196 9454 30248 9460
rect 30104 8968 30156 8974
rect 30104 8910 30156 8916
rect 30116 8634 30144 8910
rect 30104 8628 30156 8634
rect 30104 8570 30156 8576
rect 30208 8566 30236 9454
rect 30196 8560 30248 8566
rect 30196 8502 30248 8508
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 30012 7880 30064 7886
rect 30012 7822 30064 7828
rect 30024 7546 30052 7822
rect 29644 7540 29696 7546
rect 29644 7482 29696 7488
rect 30012 7540 30064 7546
rect 30012 7482 30064 7488
rect 29276 5840 29328 5846
rect 29276 5782 29328 5788
rect 29184 5772 29236 5778
rect 29184 5714 29236 5720
rect 28448 5296 28500 5302
rect 28448 5238 28500 5244
rect 28264 5160 28316 5166
rect 28264 5102 28316 5108
rect 29196 5098 29224 5714
rect 29288 5234 29316 5782
rect 30300 5642 30328 10610
rect 30380 10124 30432 10130
rect 30576 10112 30604 12192
rect 30656 11688 30708 11694
rect 30656 11630 30708 11636
rect 30668 11354 30696 11630
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30656 11008 30708 11014
rect 30656 10950 30708 10956
rect 30432 10084 30604 10112
rect 30380 10066 30432 10072
rect 30668 10062 30696 10950
rect 30760 10266 30788 13738
rect 30748 10260 30800 10266
rect 30748 10202 30800 10208
rect 30656 10056 30708 10062
rect 30656 9998 30708 10004
rect 30840 9920 30892 9926
rect 30840 9862 30892 9868
rect 30852 9586 30880 9862
rect 30748 9580 30800 9586
rect 30748 9522 30800 9528
rect 30840 9580 30892 9586
rect 30840 9522 30892 9528
rect 30654 9480 30710 9489
rect 30654 9415 30710 9424
rect 30380 8900 30432 8906
rect 30380 8842 30432 8848
rect 30392 8072 30420 8842
rect 30392 8044 30604 8072
rect 30392 7886 30420 8044
rect 30472 7948 30524 7954
rect 30472 7890 30524 7896
rect 30380 7880 30432 7886
rect 30380 7822 30432 7828
rect 30484 6798 30512 7890
rect 30576 7750 30604 8044
rect 30564 7744 30616 7750
rect 30564 7686 30616 7692
rect 30576 6798 30604 7686
rect 30668 7410 30696 9415
rect 30760 9178 30788 9522
rect 30944 9450 30972 16102
rect 31128 15026 31156 19343
rect 31312 18766 31340 25094
rect 31864 24886 31892 25434
rect 31852 24880 31904 24886
rect 31852 24822 31904 24828
rect 32600 24154 32628 31726
rect 32784 30802 32812 34478
rect 33152 33658 33180 35974
rect 33508 35692 33560 35698
rect 33508 35634 33560 35640
rect 33324 35488 33376 35494
rect 33324 35430 33376 35436
rect 33336 35154 33364 35430
rect 33324 35148 33376 35154
rect 33324 35090 33376 35096
rect 33416 35148 33468 35154
rect 33416 35090 33468 35096
rect 33428 35018 33456 35090
rect 33416 35012 33468 35018
rect 33416 34954 33468 34960
rect 33324 34944 33376 34950
rect 33324 34886 33376 34892
rect 33336 34746 33364 34886
rect 33520 34746 33548 35634
rect 33704 35154 33732 36722
rect 34060 36576 34112 36582
rect 34060 36518 34112 36524
rect 34072 36378 34100 36518
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34060 36372 34112 36378
rect 34060 36314 34112 36320
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 33692 35148 33744 35154
rect 33692 35090 33744 35096
rect 33324 34740 33376 34746
rect 33324 34682 33376 34688
rect 33508 34740 33560 34746
rect 33508 34682 33560 34688
rect 36912 34604 36964 34610
rect 36912 34546 36964 34552
rect 34152 34536 34204 34542
rect 34152 34478 34204 34484
rect 33876 33992 33928 33998
rect 33876 33934 33928 33940
rect 33324 33856 33376 33862
rect 33324 33798 33376 33804
rect 33140 33652 33192 33658
rect 33140 33594 33192 33600
rect 33336 33522 33364 33798
rect 33888 33658 33916 33934
rect 34164 33658 34192 34478
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34336 33992 34388 33998
rect 34336 33934 34388 33940
rect 33876 33652 33928 33658
rect 33876 33594 33928 33600
rect 34152 33652 34204 33658
rect 34152 33594 34204 33600
rect 33324 33516 33376 33522
rect 33324 33458 33376 33464
rect 34244 33516 34296 33522
rect 34244 33458 34296 33464
rect 34060 33448 34112 33454
rect 34060 33390 34112 33396
rect 33232 33312 33284 33318
rect 33232 33254 33284 33260
rect 32956 32904 33008 32910
rect 32956 32846 33008 32852
rect 32864 32292 32916 32298
rect 32864 32234 32916 32240
rect 32772 30796 32824 30802
rect 32772 30738 32824 30744
rect 32680 27396 32732 27402
rect 32680 27338 32732 27344
rect 32692 26382 32720 27338
rect 32680 26376 32732 26382
rect 32680 26318 32732 26324
rect 32772 26308 32824 26314
rect 32772 26250 32824 26256
rect 32680 26240 32732 26246
rect 32680 26182 32732 26188
rect 32692 25838 32720 26182
rect 32784 25906 32812 26250
rect 32772 25900 32824 25906
rect 32772 25842 32824 25848
rect 32680 25832 32732 25838
rect 32680 25774 32732 25780
rect 32508 24126 32628 24154
rect 32772 24200 32824 24206
rect 32772 24142 32824 24148
rect 31484 24064 31536 24070
rect 31484 24006 31536 24012
rect 32404 24064 32456 24070
rect 32404 24006 32456 24012
rect 31496 23866 31524 24006
rect 31484 23860 31536 23866
rect 31484 23802 31536 23808
rect 32036 23316 32088 23322
rect 32036 23258 32088 23264
rect 31852 22976 31904 22982
rect 31852 22918 31904 22924
rect 31864 22574 31892 22918
rect 31852 22568 31904 22574
rect 31852 22510 31904 22516
rect 31864 22030 31892 22510
rect 31944 22160 31996 22166
rect 31944 22102 31996 22108
rect 31852 22024 31904 22030
rect 31852 21966 31904 21972
rect 31956 21554 31984 22102
rect 32048 22030 32076 23258
rect 32416 23118 32444 24006
rect 32508 23225 32536 24126
rect 32588 24064 32640 24070
rect 32640 24024 32720 24052
rect 32588 24006 32640 24012
rect 32494 23216 32550 23225
rect 32494 23151 32550 23160
rect 32404 23112 32456 23118
rect 32404 23054 32456 23060
rect 32496 23112 32548 23118
rect 32496 23054 32548 23060
rect 32416 22642 32444 23054
rect 32508 22778 32536 23054
rect 32588 22976 32640 22982
rect 32588 22918 32640 22924
rect 32496 22772 32548 22778
rect 32496 22714 32548 22720
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 32404 22636 32456 22642
rect 32404 22578 32456 22584
rect 32036 22024 32088 22030
rect 32036 21966 32088 21972
rect 31944 21548 31996 21554
rect 31944 21490 31996 21496
rect 32036 20528 32088 20534
rect 32036 20470 32088 20476
rect 32048 20058 32076 20470
rect 32036 20052 32088 20058
rect 32036 19994 32088 20000
rect 31576 19848 31628 19854
rect 31576 19790 31628 19796
rect 31300 18760 31352 18766
rect 31300 18702 31352 18708
rect 31392 18760 31444 18766
rect 31392 18702 31444 18708
rect 31208 18624 31260 18630
rect 31208 18566 31260 18572
rect 31220 18426 31248 18566
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31312 18358 31340 18702
rect 31300 18352 31352 18358
rect 31300 18294 31352 18300
rect 31208 17876 31260 17882
rect 31208 17818 31260 17824
rect 31220 16794 31248 17818
rect 31312 17746 31340 18294
rect 31404 17882 31432 18702
rect 31588 18222 31616 19790
rect 32036 18284 32088 18290
rect 32036 18226 32088 18232
rect 31576 18216 31628 18222
rect 31576 18158 31628 18164
rect 31392 17876 31444 17882
rect 31392 17818 31444 17824
rect 31300 17740 31352 17746
rect 31300 17682 31352 17688
rect 31208 16788 31260 16794
rect 31208 16730 31260 16736
rect 31484 16584 31536 16590
rect 31484 16526 31536 16532
rect 31392 15904 31444 15910
rect 31392 15846 31444 15852
rect 31404 15706 31432 15846
rect 31392 15700 31444 15706
rect 31392 15642 31444 15648
rect 31116 15020 31168 15026
rect 31116 14962 31168 14968
rect 31024 14816 31076 14822
rect 31024 14758 31076 14764
rect 31036 14550 31064 14758
rect 31024 14544 31076 14550
rect 31024 14486 31076 14492
rect 30932 9444 30984 9450
rect 30932 9386 30984 9392
rect 30748 9172 30800 9178
rect 30748 9114 30800 9120
rect 30932 8832 30984 8838
rect 30932 8774 30984 8780
rect 30840 8084 30892 8090
rect 30840 8026 30892 8032
rect 30852 7886 30880 8026
rect 30944 7886 30972 8774
rect 31024 8424 31076 8430
rect 31024 8366 31076 8372
rect 31036 7886 31064 8366
rect 31128 7954 31156 14962
rect 31392 14816 31444 14822
rect 31392 14758 31444 14764
rect 31404 14278 31432 14758
rect 31208 14272 31260 14278
rect 31208 14214 31260 14220
rect 31392 14272 31444 14278
rect 31392 14214 31444 14220
rect 31220 13462 31248 14214
rect 31496 14074 31524 16526
rect 31588 14550 31616 18158
rect 31760 18080 31812 18086
rect 31760 18022 31812 18028
rect 31772 16998 31800 18022
rect 32048 17678 32076 18226
rect 32140 18154 32168 22578
rect 32600 22438 32628 22918
rect 32496 22432 32548 22438
rect 32496 22374 32548 22380
rect 32588 22432 32640 22438
rect 32588 22374 32640 22380
rect 32508 21842 32536 22374
rect 32600 21962 32628 22374
rect 32692 22030 32720 24024
rect 32784 22166 32812 24142
rect 32772 22160 32824 22166
rect 32772 22102 32824 22108
rect 32876 22094 32904 32234
rect 32968 31142 32996 32846
rect 33244 32434 33272 33254
rect 33324 33108 33376 33114
rect 33324 33050 33376 33056
rect 33140 32428 33192 32434
rect 33140 32370 33192 32376
rect 33232 32428 33284 32434
rect 33232 32370 33284 32376
rect 32956 31136 33008 31142
rect 32956 31078 33008 31084
rect 32968 30394 32996 31078
rect 33152 30954 33180 32370
rect 33060 30926 33180 30954
rect 33336 30938 33364 33050
rect 33782 32464 33838 32473
rect 33782 32399 33838 32408
rect 33324 30932 33376 30938
rect 32956 30388 33008 30394
rect 32956 30330 33008 30336
rect 33060 30326 33088 30926
rect 33324 30874 33376 30880
rect 33140 30796 33192 30802
rect 33140 30738 33192 30744
rect 33048 30320 33100 30326
rect 33048 30262 33100 30268
rect 32956 30048 33008 30054
rect 32956 29990 33008 29996
rect 32968 24834 32996 29990
rect 33048 29164 33100 29170
rect 33048 29106 33100 29112
rect 33060 28218 33088 29106
rect 33048 28212 33100 28218
rect 33048 28154 33100 28160
rect 33152 28014 33180 30738
rect 33692 30660 33744 30666
rect 33692 30602 33744 30608
rect 33324 30592 33376 30598
rect 33324 30534 33376 30540
rect 33232 30320 33284 30326
rect 33232 30262 33284 30268
rect 33244 29102 33272 30262
rect 33336 30122 33364 30534
rect 33324 30116 33376 30122
rect 33324 30058 33376 30064
rect 33336 29510 33364 30058
rect 33704 29617 33732 30602
rect 33690 29608 33746 29617
rect 33690 29543 33746 29552
rect 33324 29504 33376 29510
rect 33324 29446 33376 29452
rect 33232 29096 33284 29102
rect 33232 29038 33284 29044
rect 33324 28620 33376 28626
rect 33324 28562 33376 28568
rect 33140 28008 33192 28014
rect 33140 27950 33192 27956
rect 33140 26988 33192 26994
rect 33140 26930 33192 26936
rect 33152 26586 33180 26930
rect 33140 26580 33192 26586
rect 33140 26522 33192 26528
rect 33336 26246 33364 28562
rect 33796 27606 33824 32399
rect 34072 30841 34100 33390
rect 34256 33318 34284 33458
rect 34244 33312 34296 33318
rect 34244 33254 34296 33260
rect 34348 32910 34376 33934
rect 36268 33924 36320 33930
rect 36268 33866 36320 33872
rect 35992 33856 36044 33862
rect 35992 33798 36044 33804
rect 34796 33312 34848 33318
rect 34796 33254 34848 33260
rect 34808 33114 34836 33254
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34796 33108 34848 33114
rect 34796 33050 34848 33056
rect 36004 32910 36032 33798
rect 36280 33522 36308 33866
rect 36924 33658 36952 34546
rect 37924 34536 37976 34542
rect 37924 34478 37976 34484
rect 37936 34105 37964 34478
rect 37922 34096 37978 34105
rect 37922 34031 37978 34040
rect 36912 33652 36964 33658
rect 36912 33594 36964 33600
rect 36268 33516 36320 33522
rect 36268 33458 36320 33464
rect 36728 33516 36780 33522
rect 36728 33458 36780 33464
rect 34336 32904 34388 32910
rect 34336 32846 34388 32852
rect 35992 32904 36044 32910
rect 35992 32846 36044 32852
rect 35624 32768 35676 32774
rect 35624 32710 35676 32716
rect 34612 32496 34664 32502
rect 34612 32438 34664 32444
rect 34624 31822 34652 32438
rect 35636 32434 35664 32710
rect 35624 32428 35676 32434
rect 35624 32370 35676 32376
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34612 31816 34664 31822
rect 34612 31758 34664 31764
rect 35440 31816 35492 31822
rect 35440 31758 35492 31764
rect 34520 31748 34572 31754
rect 34520 31690 34572 31696
rect 34532 31346 34560 31690
rect 34520 31340 34572 31346
rect 34520 31282 34572 31288
rect 34152 31272 34204 31278
rect 34152 31214 34204 31220
rect 34164 30938 34192 31214
rect 34152 30932 34204 30938
rect 34152 30874 34204 30880
rect 34058 30832 34114 30841
rect 33968 30796 34020 30802
rect 34058 30767 34114 30776
rect 33968 30738 34020 30744
rect 33980 28626 34008 30738
rect 34072 29782 34100 30767
rect 34060 29776 34112 29782
rect 34060 29718 34112 29724
rect 34244 29776 34296 29782
rect 34244 29718 34296 29724
rect 33968 28620 34020 28626
rect 33968 28562 34020 28568
rect 34060 28484 34112 28490
rect 34060 28426 34112 28432
rect 33876 28008 33928 28014
rect 33876 27950 33928 27956
rect 33784 27600 33836 27606
rect 33784 27542 33836 27548
rect 33600 27328 33652 27334
rect 33600 27270 33652 27276
rect 33612 27062 33640 27270
rect 33600 27056 33652 27062
rect 33600 26998 33652 27004
rect 33784 26920 33836 26926
rect 33784 26862 33836 26868
rect 33796 26382 33824 26862
rect 33888 26450 33916 27950
rect 34072 27130 34100 28426
rect 34152 28416 34204 28422
rect 34152 28358 34204 28364
rect 34164 28082 34192 28358
rect 34152 28076 34204 28082
rect 34152 28018 34204 28024
rect 34256 27962 34284 29718
rect 34336 29572 34388 29578
rect 34336 29514 34388 29520
rect 34348 29238 34376 29514
rect 34520 29504 34572 29510
rect 34520 29446 34572 29452
rect 34336 29232 34388 29238
rect 34336 29174 34388 29180
rect 34164 27934 34284 27962
rect 34060 27124 34112 27130
rect 34060 27066 34112 27072
rect 33876 26444 33928 26450
rect 33876 26386 33928 26392
rect 33784 26376 33836 26382
rect 33784 26318 33836 26324
rect 33324 26240 33376 26246
rect 33324 26182 33376 26188
rect 33322 25936 33378 25945
rect 33232 25900 33284 25906
rect 33322 25871 33324 25880
rect 33232 25842 33284 25848
rect 33376 25871 33378 25880
rect 33324 25842 33376 25848
rect 33244 24954 33272 25842
rect 34164 25838 34192 27934
rect 34348 27606 34376 29174
rect 34532 29170 34560 29446
rect 34520 29164 34572 29170
rect 34520 29106 34572 29112
rect 34428 28484 34480 28490
rect 34428 28426 34480 28432
rect 34440 28218 34468 28426
rect 34520 28416 34572 28422
rect 34520 28358 34572 28364
rect 34428 28212 34480 28218
rect 34428 28154 34480 28160
rect 34532 28082 34560 28358
rect 34624 28218 34652 31758
rect 34796 31680 34848 31686
rect 34796 31622 34848 31628
rect 35256 31680 35308 31686
rect 35256 31622 35308 31628
rect 34808 31482 34836 31622
rect 34796 31476 34848 31482
rect 34796 31418 34848 31424
rect 35268 31278 35296 31622
rect 35256 31272 35308 31278
rect 35256 31214 35308 31220
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35452 30938 35480 31758
rect 35992 31136 36044 31142
rect 35992 31078 36044 31084
rect 35440 30932 35492 30938
rect 35440 30874 35492 30880
rect 36004 30326 36032 31078
rect 35992 30320 36044 30326
rect 35992 30262 36044 30268
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34796 29640 34848 29646
rect 34796 29582 34848 29588
rect 34808 29306 34836 29582
rect 34980 29572 35032 29578
rect 34980 29514 35032 29520
rect 34796 29300 34848 29306
rect 34796 29242 34848 29248
rect 34992 29170 35020 29514
rect 36004 29510 36032 30262
rect 36280 29753 36308 33458
rect 36740 32570 36768 33458
rect 36728 32564 36780 32570
rect 36728 32506 36780 32512
rect 36544 31272 36596 31278
rect 36544 31214 36596 31220
rect 36556 30666 36584 31214
rect 36544 30660 36596 30666
rect 36544 30602 36596 30608
rect 36266 29744 36322 29753
rect 36266 29679 36322 29688
rect 36634 29744 36690 29753
rect 36634 29679 36690 29688
rect 35992 29504 36044 29510
rect 35992 29446 36044 29452
rect 34980 29164 35032 29170
rect 34980 29106 35032 29112
rect 34704 29028 34756 29034
rect 34704 28970 34756 28976
rect 34716 28642 34744 28970
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34716 28614 34836 28642
rect 34704 28552 34756 28558
rect 34704 28494 34756 28500
rect 34716 28218 34744 28494
rect 34612 28212 34664 28218
rect 34612 28154 34664 28160
rect 34704 28212 34756 28218
rect 34704 28154 34756 28160
rect 34520 28076 34572 28082
rect 34520 28018 34572 28024
rect 34624 27674 34652 28154
rect 34612 27668 34664 27674
rect 34612 27610 34664 27616
rect 34336 27600 34388 27606
rect 34336 27542 34388 27548
rect 34244 26308 34296 26314
rect 34244 26250 34296 26256
rect 34256 25838 34284 26250
rect 34348 26042 34376 27542
rect 34704 26376 34756 26382
rect 34704 26318 34756 26324
rect 34716 26042 34744 26318
rect 34336 26036 34388 26042
rect 34336 25978 34388 25984
rect 34704 26036 34756 26042
rect 34704 25978 34756 25984
rect 34808 25922 34836 28614
rect 36004 28490 36032 29446
rect 36648 29170 36676 29679
rect 36636 29164 36688 29170
rect 36636 29106 36688 29112
rect 36820 29164 36872 29170
rect 36820 29106 36872 29112
rect 35992 28484 36044 28490
rect 35992 28426 36044 28432
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 36004 26994 36032 28426
rect 35992 26988 36044 26994
rect 35992 26930 36044 26936
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34980 26376 35032 26382
rect 34980 26318 35032 26324
rect 34992 26042 35020 26318
rect 36004 26314 36032 26930
rect 35992 26308 36044 26314
rect 35992 26250 36044 26256
rect 36636 26308 36688 26314
rect 36636 26250 36688 26256
rect 34980 26036 35032 26042
rect 34980 25978 35032 25984
rect 34624 25894 34836 25922
rect 34152 25832 34204 25838
rect 34152 25774 34204 25780
rect 34244 25832 34296 25838
rect 34244 25774 34296 25780
rect 33324 25492 33376 25498
rect 33324 25434 33376 25440
rect 33336 24954 33364 25434
rect 33232 24948 33284 24954
rect 33232 24890 33284 24896
rect 33324 24948 33376 24954
rect 33324 24890 33376 24896
rect 32968 24806 33180 24834
rect 33152 24750 33180 24806
rect 33784 24812 33836 24818
rect 33784 24754 33836 24760
rect 33048 24744 33100 24750
rect 33048 24686 33100 24692
rect 33140 24744 33192 24750
rect 33324 24744 33376 24750
rect 33140 24686 33192 24692
rect 33244 24704 33324 24732
rect 33060 24274 33088 24686
rect 33244 24392 33272 24704
rect 33324 24686 33376 24692
rect 33324 24608 33376 24614
rect 33324 24550 33376 24556
rect 33416 24608 33468 24614
rect 33416 24550 33468 24556
rect 33152 24364 33272 24392
rect 33048 24268 33100 24274
rect 33048 24210 33100 24216
rect 32956 24200 33008 24206
rect 32956 24142 33008 24148
rect 32968 23866 32996 24142
rect 32956 23860 33008 23866
rect 32956 23802 33008 23808
rect 32968 23118 32996 23802
rect 33060 23594 33088 24210
rect 33152 24206 33180 24364
rect 33336 24206 33364 24550
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 33140 24064 33192 24070
rect 33140 24006 33192 24012
rect 33152 23866 33180 24006
rect 33140 23860 33192 23866
rect 33140 23802 33192 23808
rect 33428 23662 33456 24550
rect 33508 24336 33560 24342
rect 33508 24278 33560 24284
rect 33416 23656 33468 23662
rect 33416 23598 33468 23604
rect 33048 23588 33100 23594
rect 33048 23530 33100 23536
rect 33232 23520 33284 23526
rect 33232 23462 33284 23468
rect 33048 23316 33100 23322
rect 33048 23258 33100 23264
rect 32956 23112 33008 23118
rect 32956 23054 33008 23060
rect 33060 22778 33088 23258
rect 33048 22772 33100 22778
rect 33048 22714 33100 22720
rect 33060 22642 33088 22714
rect 33244 22642 33272 23462
rect 33324 23044 33376 23050
rect 33324 22986 33376 22992
rect 33336 22642 33364 22986
rect 33048 22636 33100 22642
rect 33048 22578 33100 22584
rect 33232 22636 33284 22642
rect 33232 22578 33284 22584
rect 33324 22636 33376 22642
rect 33324 22578 33376 22584
rect 32956 22568 33008 22574
rect 32956 22510 33008 22516
rect 32968 22250 32996 22510
rect 33232 22500 33284 22506
rect 33232 22442 33284 22448
rect 32968 22222 33088 22250
rect 33244 22234 33272 22442
rect 33336 22234 33364 22578
rect 32876 22066 32996 22094
rect 32680 22024 32732 22030
rect 32680 21966 32732 21972
rect 32588 21956 32640 21962
rect 32588 21898 32640 21904
rect 32508 21814 32720 21842
rect 32588 21684 32640 21690
rect 32588 21626 32640 21632
rect 32312 21004 32364 21010
rect 32312 20946 32364 20952
rect 32324 18630 32352 20946
rect 32600 20466 32628 21626
rect 32692 21554 32720 21814
rect 32680 21548 32732 21554
rect 32680 21490 32732 21496
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 32968 19922 32996 22066
rect 33060 21010 33088 22222
rect 33232 22228 33284 22234
rect 33232 22170 33284 22176
rect 33324 22228 33376 22234
rect 33324 22170 33376 22176
rect 33244 22098 33272 22170
rect 33232 22092 33284 22098
rect 33232 22034 33284 22040
rect 33336 21554 33364 22170
rect 33520 22098 33548 24278
rect 33796 24206 33824 24754
rect 34164 24614 34192 25774
rect 34336 25288 34388 25294
rect 34336 25230 34388 25236
rect 34348 24954 34376 25230
rect 34336 24948 34388 24954
rect 34336 24890 34388 24896
rect 34152 24608 34204 24614
rect 34152 24550 34204 24556
rect 33784 24200 33836 24206
rect 33784 24142 33836 24148
rect 34624 23730 34652 25894
rect 34704 25764 34756 25770
rect 34704 25706 34756 25712
rect 34716 25430 34744 25706
rect 34796 25696 34848 25702
rect 34796 25638 34848 25644
rect 34704 25424 34756 25430
rect 34704 25366 34756 25372
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34624 23322 34652 23666
rect 34612 23316 34664 23322
rect 34612 23258 34664 23264
rect 34808 23202 34836 25638
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36004 25226 36032 26250
rect 36648 25906 36676 26250
rect 36636 25900 36688 25906
rect 36636 25842 36688 25848
rect 35992 25220 36044 25226
rect 35992 25162 36044 25168
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35348 23656 35400 23662
rect 35348 23598 35400 23604
rect 35808 23656 35860 23662
rect 35808 23598 35860 23604
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34808 23174 35112 23202
rect 35084 23118 35112 23174
rect 34980 23112 35032 23118
rect 34980 23054 35032 23060
rect 35072 23112 35124 23118
rect 35072 23054 35124 23060
rect 34336 22976 34388 22982
rect 34336 22918 34388 22924
rect 33508 22092 33560 22098
rect 33508 22034 33560 22040
rect 33784 21684 33836 21690
rect 33784 21626 33836 21632
rect 33796 21554 33824 21626
rect 33324 21548 33376 21554
rect 33324 21490 33376 21496
rect 33600 21548 33652 21554
rect 33600 21490 33652 21496
rect 33784 21548 33836 21554
rect 33784 21490 33836 21496
rect 33612 21434 33640 21490
rect 33520 21406 33640 21434
rect 33232 21344 33284 21350
rect 33232 21286 33284 21292
rect 33048 21004 33100 21010
rect 33048 20946 33100 20952
rect 33244 20398 33272 21286
rect 33520 21146 33548 21406
rect 33508 21140 33560 21146
rect 33508 21082 33560 21088
rect 33416 20936 33468 20942
rect 33416 20878 33468 20884
rect 33324 20868 33376 20874
rect 33324 20810 33376 20816
rect 33336 20534 33364 20810
rect 33324 20528 33376 20534
rect 33324 20470 33376 20476
rect 33232 20392 33284 20398
rect 33232 20334 33284 20340
rect 33140 20324 33192 20330
rect 33140 20266 33192 20272
rect 33152 19922 33180 20266
rect 32956 19916 33008 19922
rect 32956 19858 33008 19864
rect 33140 19916 33192 19922
rect 33140 19858 33192 19864
rect 32968 19514 32996 19858
rect 32956 19508 33008 19514
rect 32956 19450 33008 19456
rect 33152 19378 33180 19858
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 33140 19168 33192 19174
rect 33140 19110 33192 19116
rect 32864 18964 32916 18970
rect 32864 18906 32916 18912
rect 32680 18760 32732 18766
rect 32680 18702 32732 18708
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32312 18624 32364 18630
rect 32312 18566 32364 18572
rect 32128 18148 32180 18154
rect 32128 18090 32180 18096
rect 32036 17672 32088 17678
rect 32036 17614 32088 17620
rect 31852 17536 31904 17542
rect 31852 17478 31904 17484
rect 31864 17202 31892 17478
rect 32048 17338 32076 17614
rect 32036 17332 32088 17338
rect 32036 17274 32088 17280
rect 32034 17232 32090 17241
rect 31852 17196 31904 17202
rect 32034 17167 32090 17176
rect 32128 17196 32180 17202
rect 31852 17138 31904 17144
rect 31864 16998 31892 17138
rect 32048 17066 32076 17167
rect 32128 17138 32180 17144
rect 32036 17060 32088 17066
rect 32036 17002 32088 17008
rect 31760 16992 31812 16998
rect 31760 16934 31812 16940
rect 31852 16992 31904 16998
rect 31852 16934 31904 16940
rect 31772 16590 31800 16934
rect 32140 16794 32168 17138
rect 32324 17134 32352 18566
rect 32692 18426 32720 18702
rect 32680 18420 32732 18426
rect 32680 18362 32732 18368
rect 32680 18284 32732 18290
rect 32784 18272 32812 18702
rect 32732 18244 32812 18272
rect 32680 18226 32732 18232
rect 32496 18216 32548 18222
rect 32496 18158 32548 18164
rect 32588 18216 32640 18222
rect 32588 18158 32640 18164
rect 32508 17882 32536 18158
rect 32496 17876 32548 17882
rect 32496 17818 32548 17824
rect 32600 17814 32628 18158
rect 32588 17808 32640 17814
rect 32588 17750 32640 17756
rect 32692 17626 32720 18226
rect 32772 18148 32824 18154
rect 32772 18090 32824 18096
rect 32508 17598 32720 17626
rect 32312 17128 32364 17134
rect 32312 17070 32364 17076
rect 32128 16788 32180 16794
rect 32128 16730 32180 16736
rect 31760 16584 31812 16590
rect 31760 16526 31812 16532
rect 32220 16040 32272 16046
rect 32220 15982 32272 15988
rect 32232 15706 32260 15982
rect 32220 15700 32272 15706
rect 32220 15642 32272 15648
rect 32232 15434 32260 15642
rect 32220 15428 32272 15434
rect 32220 15370 32272 15376
rect 31576 14544 31628 14550
rect 31576 14486 31628 14492
rect 31484 14068 31536 14074
rect 31484 14010 31536 14016
rect 31208 13456 31260 13462
rect 31208 13398 31260 13404
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 31220 12986 31248 13262
rect 31300 13252 31352 13258
rect 31300 13194 31352 13200
rect 31208 12980 31260 12986
rect 31208 12922 31260 12928
rect 31208 12844 31260 12850
rect 31312 12832 31340 13194
rect 31260 12804 31340 12832
rect 31392 12844 31444 12850
rect 31208 12786 31260 12792
rect 31392 12786 31444 12792
rect 31404 9586 31432 12786
rect 31588 12434 31616 14486
rect 31668 14476 31720 14482
rect 31668 14418 31720 14424
rect 31680 13258 31708 14418
rect 31852 13728 31904 13734
rect 31852 13670 31904 13676
rect 31668 13252 31720 13258
rect 31668 13194 31720 13200
rect 31680 12782 31708 13194
rect 31864 12986 31892 13670
rect 32128 13456 32180 13462
rect 32128 13398 32180 13404
rect 31852 12980 31904 12986
rect 31852 12922 31904 12928
rect 31668 12776 31720 12782
rect 31668 12718 31720 12724
rect 32036 12708 32088 12714
rect 32036 12650 32088 12656
rect 31496 12406 31616 12434
rect 31760 12436 31812 12442
rect 31392 9580 31444 9586
rect 31392 9522 31444 9528
rect 31404 8634 31432 9522
rect 31392 8628 31444 8634
rect 31392 8570 31444 8576
rect 31496 8090 31524 12406
rect 31760 12378 31812 12384
rect 31772 11286 31800 12378
rect 31760 11280 31812 11286
rect 31760 11222 31812 11228
rect 31852 11144 31904 11150
rect 31852 11086 31904 11092
rect 31864 10674 31892 11086
rect 31852 10668 31904 10674
rect 31852 10610 31904 10616
rect 31576 9376 31628 9382
rect 31576 9318 31628 9324
rect 31668 9376 31720 9382
rect 31668 9318 31720 9324
rect 31588 9178 31616 9318
rect 31576 9172 31628 9178
rect 31576 9114 31628 9120
rect 31680 9058 31708 9318
rect 31588 9030 31708 9058
rect 31484 8084 31536 8090
rect 31484 8026 31536 8032
rect 31116 7948 31168 7954
rect 31116 7890 31168 7896
rect 30840 7880 30892 7886
rect 30840 7822 30892 7828
rect 30932 7880 30984 7886
rect 30932 7822 30984 7828
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 30656 7404 30708 7410
rect 30656 7346 30708 7352
rect 30852 6798 30880 7822
rect 30944 7002 30972 7822
rect 30932 6996 30984 7002
rect 30932 6938 30984 6944
rect 30472 6792 30524 6798
rect 30472 6734 30524 6740
rect 30564 6792 30616 6798
rect 30564 6734 30616 6740
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30484 5914 30512 6734
rect 31036 6458 31064 7822
rect 31208 7744 31260 7750
rect 31208 7686 31260 7692
rect 31220 7546 31248 7686
rect 31208 7540 31260 7546
rect 31208 7482 31260 7488
rect 31588 7478 31616 9030
rect 31864 8974 31892 10610
rect 32048 10554 32076 12650
rect 32140 11354 32168 13398
rect 32324 12306 32352 17070
rect 32508 16522 32536 17598
rect 32588 17128 32640 17134
rect 32588 17070 32640 17076
rect 32600 16794 32628 17070
rect 32588 16788 32640 16794
rect 32588 16730 32640 16736
rect 32588 16652 32640 16658
rect 32588 16594 32640 16600
rect 32496 16516 32548 16522
rect 32496 16458 32548 16464
rect 32404 13864 32456 13870
rect 32404 13806 32456 13812
rect 32416 13530 32444 13806
rect 32404 13524 32456 13530
rect 32404 13466 32456 13472
rect 32508 12442 32536 16458
rect 32600 15706 32628 16594
rect 32588 15700 32640 15706
rect 32640 15660 32720 15688
rect 32588 15642 32640 15648
rect 32588 15360 32640 15366
rect 32588 15302 32640 15308
rect 32600 15162 32628 15302
rect 32588 15156 32640 15162
rect 32588 15098 32640 15104
rect 32588 13728 32640 13734
rect 32588 13670 32640 13676
rect 32600 13258 32628 13670
rect 32588 13252 32640 13258
rect 32588 13194 32640 13200
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 32312 12300 32364 12306
rect 32312 12242 32364 12248
rect 32600 12102 32628 13194
rect 32692 12782 32720 15660
rect 32680 12776 32732 12782
rect 32680 12718 32732 12724
rect 32680 12436 32732 12442
rect 32680 12378 32732 12384
rect 32588 12096 32640 12102
rect 32588 12038 32640 12044
rect 32692 11898 32720 12378
rect 32784 12322 32812 18090
rect 32876 17338 32904 18906
rect 33152 18834 33180 19110
rect 33140 18828 33192 18834
rect 33140 18770 33192 18776
rect 32956 18760 33008 18766
rect 32956 18702 33008 18708
rect 32968 18630 32996 18702
rect 32956 18624 33008 18630
rect 32956 18566 33008 18572
rect 33140 18624 33192 18630
rect 33140 18566 33192 18572
rect 33152 18358 33180 18566
rect 33140 18352 33192 18358
rect 33140 18294 33192 18300
rect 33428 17678 33456 20878
rect 33520 19334 33548 21082
rect 34348 21078 34376 22918
rect 34992 22642 35020 23054
rect 35084 22778 35112 23054
rect 35072 22772 35124 22778
rect 35072 22714 35124 22720
rect 35360 22642 35388 23598
rect 35820 23186 35848 23598
rect 35808 23180 35860 23186
rect 35808 23122 35860 23128
rect 36084 22976 36136 22982
rect 36084 22918 36136 22924
rect 36176 22976 36228 22982
rect 36176 22918 36228 22924
rect 34428 22636 34480 22642
rect 34428 22578 34480 22584
rect 34980 22636 35032 22642
rect 34980 22578 35032 22584
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 35808 22636 35860 22642
rect 35808 22578 35860 22584
rect 34440 22030 34468 22578
rect 34796 22432 34848 22438
rect 34796 22374 34848 22380
rect 34808 22030 34836 22374
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34428 22024 34480 22030
rect 34428 21966 34480 21972
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 35256 22024 35308 22030
rect 35256 21966 35308 21972
rect 34704 21888 34756 21894
rect 34704 21830 34756 21836
rect 34610 21720 34666 21729
rect 34716 21690 34744 21830
rect 35268 21690 35296 21966
rect 34610 21655 34666 21664
rect 34704 21684 34756 21690
rect 34336 21072 34388 21078
rect 34336 21014 34388 21020
rect 34428 20392 34480 20398
rect 34428 20334 34480 20340
rect 34152 19372 34204 19378
rect 33520 19306 33824 19334
rect 34152 19314 34204 19320
rect 33796 18329 33824 19306
rect 33968 18760 34020 18766
rect 33968 18702 34020 18708
rect 33782 18320 33838 18329
rect 33782 18255 33838 18264
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 32864 17332 32916 17338
rect 32864 17274 32916 17280
rect 33048 17332 33100 17338
rect 33048 17274 33100 17280
rect 32862 17232 32918 17241
rect 32862 17167 32864 17176
rect 32916 17167 32918 17176
rect 32864 17138 32916 17144
rect 32864 15700 32916 15706
rect 32864 15642 32916 15648
rect 32876 15502 32904 15642
rect 32864 15496 32916 15502
rect 32864 15438 32916 15444
rect 32876 14074 32904 15438
rect 33060 15026 33088 17274
rect 33428 16998 33456 17614
rect 33796 17542 33824 18255
rect 33980 18086 34008 18702
rect 34164 18426 34192 19314
rect 34440 19242 34468 20334
rect 34520 20324 34572 20330
rect 34520 20266 34572 20272
rect 34428 19236 34480 19242
rect 34428 19178 34480 19184
rect 34440 18970 34468 19178
rect 34428 18964 34480 18970
rect 34428 18906 34480 18912
rect 34152 18420 34204 18426
rect 34152 18362 34204 18368
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 33980 17678 34008 18022
rect 34060 17808 34112 17814
rect 34060 17750 34112 17756
rect 33968 17672 34020 17678
rect 33968 17614 34020 17620
rect 33784 17536 33836 17542
rect 33784 17478 33836 17484
rect 33796 17270 33824 17478
rect 33980 17338 34008 17614
rect 33968 17332 34020 17338
rect 33968 17274 34020 17280
rect 33784 17264 33836 17270
rect 33784 17206 33836 17212
rect 33416 16992 33468 16998
rect 33416 16934 33468 16940
rect 33416 15496 33468 15502
rect 33416 15438 33468 15444
rect 33048 15020 33100 15026
rect 33048 14962 33100 14968
rect 32956 14952 33008 14958
rect 32956 14894 33008 14900
rect 32968 14618 32996 14894
rect 32956 14612 33008 14618
rect 32956 14554 33008 14560
rect 32864 14068 32916 14074
rect 32864 14010 32916 14016
rect 32956 13932 33008 13938
rect 32956 13874 33008 13880
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 32864 13320 32916 13326
rect 32864 13262 32916 13268
rect 32876 12986 32904 13262
rect 32968 13190 32996 13874
rect 33140 13728 33192 13734
rect 33140 13670 33192 13676
rect 33152 13326 33180 13670
rect 33244 13530 33272 13874
rect 33428 13530 33456 15438
rect 33796 14278 33824 17206
rect 34072 17134 34100 17750
rect 34532 17270 34560 20266
rect 34624 20074 34652 21655
rect 34704 21626 34756 21632
rect 35256 21684 35308 21690
rect 35256 21626 35308 21632
rect 35360 21622 35388 22578
rect 35624 22092 35676 22098
rect 35624 22034 35676 22040
rect 35348 21616 35400 21622
rect 35348 21558 35400 21564
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35256 21140 35308 21146
rect 35256 21082 35308 21088
rect 35268 20942 35296 21082
rect 35360 21078 35388 21558
rect 35636 21486 35664 22034
rect 35716 21888 35768 21894
rect 35716 21830 35768 21836
rect 35728 21554 35756 21830
rect 35820 21554 35848 22578
rect 35900 22432 35952 22438
rect 35900 22374 35952 22380
rect 35716 21548 35768 21554
rect 35716 21490 35768 21496
rect 35808 21548 35860 21554
rect 35808 21490 35860 21496
rect 35624 21480 35676 21486
rect 35624 21422 35676 21428
rect 35440 21344 35492 21350
rect 35440 21286 35492 21292
rect 35452 21146 35480 21286
rect 35440 21140 35492 21146
rect 35440 21082 35492 21088
rect 35348 21072 35400 21078
rect 35400 21020 35480 21026
rect 35348 21014 35480 21020
rect 35360 20998 35480 21014
rect 35452 20942 35480 20998
rect 35256 20936 35308 20942
rect 35256 20878 35308 20884
rect 35440 20936 35492 20942
rect 35440 20878 35492 20884
rect 34796 20256 34848 20262
rect 34796 20198 34848 20204
rect 34624 20058 34744 20074
rect 34624 20052 34756 20058
rect 34624 20046 34704 20052
rect 34704 19994 34756 20000
rect 34612 19984 34664 19990
rect 34612 19926 34664 19932
rect 34520 17264 34572 17270
rect 34520 17206 34572 17212
rect 34532 17134 34560 17206
rect 34060 17128 34112 17134
rect 34060 17070 34112 17076
rect 34520 17128 34572 17134
rect 34520 17070 34572 17076
rect 34520 16516 34572 16522
rect 34520 16458 34572 16464
rect 34532 15910 34560 16458
rect 34520 15904 34572 15910
rect 34520 15846 34572 15852
rect 34624 15502 34652 19926
rect 34716 15502 34744 19994
rect 34808 19718 34836 20198
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35164 20052 35216 20058
rect 35164 19994 35216 20000
rect 35176 19854 35204 19994
rect 35636 19922 35664 21422
rect 35728 20058 35756 21490
rect 35820 20602 35848 21490
rect 35808 20596 35860 20602
rect 35808 20538 35860 20544
rect 35912 20466 35940 22374
rect 36096 22098 36124 22918
rect 36188 22710 36216 22918
rect 36452 22772 36504 22778
rect 36280 22732 36452 22760
rect 36176 22704 36228 22710
rect 36176 22646 36228 22652
rect 36280 22642 36308 22732
rect 36452 22714 36504 22720
rect 36268 22636 36320 22642
rect 36268 22578 36320 22584
rect 36452 22432 36504 22438
rect 36452 22374 36504 22380
rect 36176 22228 36228 22234
rect 36176 22170 36228 22176
rect 36084 22092 36136 22098
rect 36084 22034 36136 22040
rect 36188 21554 36216 22170
rect 36464 22098 36492 22374
rect 36452 22092 36504 22098
rect 36452 22034 36504 22040
rect 36464 21554 36492 22034
rect 36176 21548 36228 21554
rect 36176 21490 36228 21496
rect 36452 21548 36504 21554
rect 36452 21490 36504 21496
rect 35900 20460 35952 20466
rect 35900 20402 35952 20408
rect 35808 20392 35860 20398
rect 35808 20334 35860 20340
rect 35820 20058 35848 20334
rect 35716 20052 35768 20058
rect 35716 19994 35768 20000
rect 35808 20052 35860 20058
rect 35808 19994 35860 20000
rect 35624 19916 35676 19922
rect 35624 19858 35676 19864
rect 35164 19848 35216 19854
rect 35164 19790 35216 19796
rect 35440 19848 35492 19854
rect 35440 19790 35492 19796
rect 34796 19712 34848 19718
rect 34796 19654 34848 19660
rect 34808 19514 34836 19654
rect 34796 19508 34848 19514
rect 34796 19450 34848 19456
rect 34796 19304 34848 19310
rect 34796 19246 34848 19252
rect 34808 18850 34836 19246
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34808 18822 35020 18850
rect 35452 18834 35480 19790
rect 34992 18630 35020 18822
rect 35440 18828 35492 18834
rect 35440 18770 35492 18776
rect 34796 18624 34848 18630
rect 34796 18566 34848 18572
rect 34980 18624 35032 18630
rect 34980 18566 35032 18572
rect 35164 18624 35216 18630
rect 35164 18566 35216 18572
rect 34808 18426 34836 18566
rect 34796 18420 34848 18426
rect 34796 18362 34848 18368
rect 34992 18290 35020 18566
rect 35176 18290 35204 18566
rect 35636 18358 35664 19858
rect 36188 19718 36216 21490
rect 35900 19712 35952 19718
rect 35900 19654 35952 19660
rect 36176 19712 36228 19718
rect 36176 19654 36228 19660
rect 35912 19514 35940 19654
rect 35900 19508 35952 19514
rect 35900 19450 35952 19456
rect 36188 19334 36216 19654
rect 36004 19306 36216 19334
rect 36648 19334 36676 25842
rect 36728 25220 36780 25226
rect 36728 25162 36780 25168
rect 36740 24886 36768 25162
rect 36728 24880 36780 24886
rect 36728 24822 36780 24828
rect 36832 21457 36860 29106
rect 37280 29028 37332 29034
rect 37280 28970 37332 28976
rect 37292 28218 37320 28970
rect 37280 28212 37332 28218
rect 37280 28154 37332 28160
rect 37556 27872 37608 27878
rect 37556 27814 37608 27820
rect 37568 22642 37596 27814
rect 37556 22636 37608 22642
rect 37556 22578 37608 22584
rect 37830 22536 37886 22545
rect 37830 22471 37832 22480
rect 37884 22471 37886 22480
rect 37832 22442 37884 22448
rect 37004 22432 37056 22438
rect 37004 22374 37056 22380
rect 37016 22094 37044 22374
rect 36924 22066 37044 22094
rect 36924 22030 36952 22066
rect 36912 22024 36964 22030
rect 36912 21966 36964 21972
rect 37188 21480 37240 21486
rect 36818 21448 36874 21457
rect 37188 21422 37240 21428
rect 36818 21383 36874 21392
rect 36648 19306 36768 19334
rect 36004 19174 36032 19306
rect 35992 19168 36044 19174
rect 35992 19110 36044 19116
rect 36740 18834 36768 19306
rect 36728 18828 36780 18834
rect 36728 18770 36780 18776
rect 36832 18698 36860 21383
rect 36820 18692 36872 18698
rect 36820 18634 36872 18640
rect 35624 18352 35676 18358
rect 35624 18294 35676 18300
rect 34980 18284 35032 18290
rect 34980 18226 35032 18232
rect 35164 18284 35216 18290
rect 35164 18226 35216 18232
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34796 16992 34848 16998
rect 34796 16934 34848 16940
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 34808 16522 34836 16934
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35360 16810 35388 16934
rect 35268 16794 35388 16810
rect 35256 16788 35388 16794
rect 35308 16782 35388 16788
rect 35440 16788 35492 16794
rect 35256 16730 35308 16736
rect 35440 16730 35492 16736
rect 34796 16516 34848 16522
rect 34796 16458 34848 16464
rect 34808 16250 34836 16458
rect 35164 16448 35216 16454
rect 35164 16390 35216 16396
rect 34796 16244 34848 16250
rect 34796 16186 34848 16192
rect 35176 16114 35204 16390
rect 35268 16250 35296 16730
rect 35256 16244 35308 16250
rect 35256 16186 35308 16192
rect 35164 16108 35216 16114
rect 35164 16050 35216 16056
rect 34796 16040 34848 16046
rect 35452 15994 35480 16730
rect 35532 16652 35584 16658
rect 35532 16594 35584 16600
rect 34796 15982 34848 15988
rect 34808 15706 34836 15982
rect 35268 15966 35480 15994
rect 35268 15910 35296 15966
rect 35256 15904 35308 15910
rect 35256 15846 35308 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35544 15706 35572 16594
rect 34796 15700 34848 15706
rect 34796 15642 34848 15648
rect 35532 15700 35584 15706
rect 35532 15642 35584 15648
rect 34796 15564 34848 15570
rect 34796 15506 34848 15512
rect 35624 15564 35676 15570
rect 35624 15506 35676 15512
rect 34612 15496 34664 15502
rect 34612 15438 34664 15444
rect 34704 15496 34756 15502
rect 34704 15438 34756 15444
rect 34808 15162 34836 15506
rect 34796 15156 34848 15162
rect 34796 15098 34848 15104
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 33784 14272 33836 14278
rect 33784 14214 33836 14220
rect 34060 14272 34112 14278
rect 34060 14214 34112 14220
rect 33508 13932 33560 13938
rect 33508 13874 33560 13880
rect 33232 13524 33284 13530
rect 33232 13466 33284 13472
rect 33416 13524 33468 13530
rect 33416 13466 33468 13472
rect 33520 13326 33548 13874
rect 33140 13320 33192 13326
rect 33140 13262 33192 13268
rect 33508 13320 33560 13326
rect 33508 13262 33560 13268
rect 33876 13320 33928 13326
rect 33876 13262 33928 13268
rect 32956 13184 33008 13190
rect 32956 13126 33008 13132
rect 32864 12980 32916 12986
rect 32864 12922 32916 12928
rect 32968 12442 32996 13126
rect 33152 12986 33180 13262
rect 33140 12980 33192 12986
rect 33140 12922 33192 12928
rect 33888 12850 33916 13262
rect 33876 12844 33928 12850
rect 33876 12786 33928 12792
rect 33324 12776 33376 12782
rect 33324 12718 33376 12724
rect 32956 12436 33008 12442
rect 32956 12378 33008 12384
rect 32784 12294 33088 12322
rect 33060 12238 33088 12294
rect 33048 12232 33100 12238
rect 33048 12174 33100 12180
rect 33232 12232 33284 12238
rect 33232 12174 33284 12180
rect 32680 11892 32732 11898
rect 32680 11834 32732 11840
rect 32220 11824 32272 11830
rect 32220 11766 32272 11772
rect 32128 11348 32180 11354
rect 32128 11290 32180 11296
rect 32232 10674 32260 11766
rect 32588 11756 32640 11762
rect 32588 11698 32640 11704
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32324 10810 32352 11086
rect 32312 10804 32364 10810
rect 32312 10746 32364 10752
rect 32220 10668 32272 10674
rect 32220 10610 32272 10616
rect 32508 10606 32536 11086
rect 32600 11014 32628 11698
rect 32692 11354 32720 11834
rect 32680 11348 32732 11354
rect 32680 11290 32732 11296
rect 32772 11144 32824 11150
rect 32772 11086 32824 11092
rect 32588 11008 32640 11014
rect 32588 10950 32640 10956
rect 32600 10810 32628 10950
rect 32588 10804 32640 10810
rect 32588 10746 32640 10752
rect 32784 10674 32812 11086
rect 32956 11008 33008 11014
rect 32956 10950 33008 10956
rect 32772 10668 32824 10674
rect 32772 10610 32824 10616
rect 32496 10600 32548 10606
rect 32048 10526 32168 10554
rect 32496 10542 32548 10548
rect 32140 10470 32168 10526
rect 32128 10464 32180 10470
rect 32128 10406 32180 10412
rect 32036 9444 32088 9450
rect 32036 9386 32088 9392
rect 32048 9042 32076 9386
rect 32036 9036 32088 9042
rect 32036 8978 32088 8984
rect 31760 8968 31812 8974
rect 31760 8910 31812 8916
rect 31852 8968 31904 8974
rect 31852 8910 31904 8916
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 31680 7818 31708 8434
rect 31772 8090 31800 8910
rect 31944 8832 31996 8838
rect 31944 8774 31996 8780
rect 31956 8566 31984 8774
rect 32048 8634 32076 8978
rect 32036 8628 32088 8634
rect 32036 8570 32088 8576
rect 31944 8560 31996 8566
rect 31944 8502 31996 8508
rect 31760 8084 31812 8090
rect 31760 8026 31812 8032
rect 31668 7812 31720 7818
rect 31668 7754 31720 7760
rect 31576 7472 31628 7478
rect 31576 7414 31628 7420
rect 31772 7410 31800 8026
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31760 7404 31812 7410
rect 31760 7346 31812 7352
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 31312 7002 31340 7278
rect 31404 7002 31432 7346
rect 31300 6996 31352 7002
rect 31300 6938 31352 6944
rect 31392 6996 31444 7002
rect 31392 6938 31444 6944
rect 31956 6882 31984 8502
rect 31772 6854 31984 6882
rect 31772 6798 31800 6854
rect 32140 6798 32168 10406
rect 32784 10266 32812 10610
rect 32864 10464 32916 10470
rect 32864 10406 32916 10412
rect 32772 10260 32824 10266
rect 32772 10202 32824 10208
rect 32784 9586 32812 10202
rect 32876 10169 32904 10406
rect 32968 10198 32996 10950
rect 32956 10192 33008 10198
rect 32862 10160 32918 10169
rect 32956 10134 33008 10140
rect 32862 10095 32918 10104
rect 32876 10062 32904 10095
rect 32864 10056 32916 10062
rect 32864 9998 32916 10004
rect 32772 9580 32824 9586
rect 32772 9522 32824 9528
rect 32772 8968 32824 8974
rect 32968 8956 32996 10134
rect 33060 9654 33088 12174
rect 33244 10606 33272 12174
rect 33232 10600 33284 10606
rect 33232 10542 33284 10548
rect 33140 9716 33192 9722
rect 33140 9658 33192 9664
rect 33048 9648 33100 9654
rect 33048 9590 33100 9596
rect 33152 9178 33180 9658
rect 33244 9382 33272 10542
rect 33232 9376 33284 9382
rect 33232 9318 33284 9324
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 33244 9058 33272 9318
rect 33336 9178 33364 12718
rect 33692 11756 33744 11762
rect 33692 11698 33744 11704
rect 33704 10810 33732 11698
rect 33692 10804 33744 10810
rect 33692 10746 33744 10752
rect 33508 10668 33560 10674
rect 33508 10610 33560 10616
rect 33520 10266 33548 10610
rect 33508 10260 33560 10266
rect 33508 10202 33560 10208
rect 34072 10062 34100 14214
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34612 11620 34664 11626
rect 34612 11562 34664 11568
rect 34624 11354 34652 11562
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34612 11348 34664 11354
rect 34612 11290 34664 11296
rect 35636 10810 35664 15506
rect 35624 10804 35676 10810
rect 35624 10746 35676 10752
rect 34428 10668 34480 10674
rect 34428 10610 34480 10616
rect 33968 10056 34020 10062
rect 33968 9998 34020 10004
rect 34060 10056 34112 10062
rect 34060 9998 34112 10004
rect 33980 9722 34008 9998
rect 33968 9716 34020 9722
rect 33968 9658 34020 9664
rect 33324 9172 33376 9178
rect 33324 9114 33376 9120
rect 33152 9030 33272 9058
rect 33152 8974 33180 9030
rect 33048 8968 33100 8974
rect 32968 8928 33048 8956
rect 32772 8910 32824 8916
rect 33048 8910 33100 8916
rect 33140 8968 33192 8974
rect 33140 8910 33192 8916
rect 32588 8356 32640 8362
rect 32588 8298 32640 8304
rect 32600 6866 32628 8298
rect 32588 6860 32640 6866
rect 32588 6802 32640 6808
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 32128 6792 32180 6798
rect 32128 6734 32180 6740
rect 31024 6452 31076 6458
rect 31024 6394 31076 6400
rect 30472 5908 30524 5914
rect 30472 5850 30524 5856
rect 31772 5710 31800 6734
rect 31944 6656 31996 6662
rect 31944 6598 31996 6604
rect 32220 6656 32272 6662
rect 32220 6598 32272 6604
rect 31760 5704 31812 5710
rect 31760 5646 31812 5652
rect 30196 5636 30248 5642
rect 30196 5578 30248 5584
rect 30288 5636 30340 5642
rect 30288 5578 30340 5584
rect 29828 5568 29880 5574
rect 29828 5510 29880 5516
rect 29840 5234 29868 5510
rect 29276 5228 29328 5234
rect 29276 5170 29328 5176
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 30104 5228 30156 5234
rect 30104 5170 30156 5176
rect 29184 5092 29236 5098
rect 29184 5034 29236 5040
rect 29196 4826 29224 5034
rect 29184 4820 29236 4826
rect 29184 4762 29236 4768
rect 29288 4690 29316 5170
rect 29828 5092 29880 5098
rect 29828 5034 29880 5040
rect 29644 5024 29696 5030
rect 29644 4966 29696 4972
rect 27988 4684 28040 4690
rect 27988 4626 28040 4632
rect 28080 4684 28132 4690
rect 28080 4626 28132 4632
rect 29276 4684 29328 4690
rect 29276 4626 29328 4632
rect 28000 4282 28028 4626
rect 29656 4622 29684 4966
rect 29840 4758 29868 5034
rect 30012 5024 30064 5030
rect 30012 4966 30064 4972
rect 30024 4826 30052 4966
rect 30012 4820 30064 4826
rect 30012 4762 30064 4768
rect 29828 4752 29880 4758
rect 29828 4694 29880 4700
rect 29644 4616 29696 4622
rect 29644 4558 29696 4564
rect 27988 4276 28040 4282
rect 27988 4218 28040 4224
rect 30116 4146 30144 5170
rect 30208 4826 30236 5578
rect 30300 5370 30328 5578
rect 30288 5364 30340 5370
rect 30288 5306 30340 5312
rect 31772 5234 31800 5646
rect 31956 5642 31984 6598
rect 32232 6322 32260 6598
rect 32220 6316 32272 6322
rect 32220 6258 32272 6264
rect 32036 6112 32088 6118
rect 32036 6054 32088 6060
rect 32048 5914 32076 6054
rect 32232 5914 32260 6258
rect 32600 6186 32628 6802
rect 32680 6792 32732 6798
rect 32680 6734 32732 6740
rect 32692 6322 32720 6734
rect 32680 6316 32732 6322
rect 32680 6258 32732 6264
rect 32784 6186 32812 8910
rect 32864 8900 32916 8906
rect 32864 8842 32916 8848
rect 32876 6866 32904 8842
rect 33060 8498 33088 8910
rect 33232 8832 33284 8838
rect 33232 8774 33284 8780
rect 33048 8492 33100 8498
rect 33048 8434 33100 8440
rect 33244 8430 33272 8774
rect 33232 8424 33284 8430
rect 33232 8366 33284 8372
rect 34072 8294 34100 9998
rect 34060 8288 34112 8294
rect 34060 8230 34112 8236
rect 33048 8016 33100 8022
rect 33048 7958 33100 7964
rect 32864 6860 32916 6866
rect 32864 6802 32916 6808
rect 33060 6798 33088 7958
rect 33140 6860 33192 6866
rect 33140 6802 33192 6808
rect 33048 6792 33100 6798
rect 33048 6734 33100 6740
rect 33152 6458 33180 6802
rect 34440 6730 34468 10610
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 36832 8906 36860 18634
rect 37096 18624 37148 18630
rect 37096 18566 37148 18572
rect 37108 18426 37136 18566
rect 37096 18420 37148 18426
rect 37096 18362 37148 18368
rect 37200 18358 37228 21422
rect 38384 20732 38436 20738
rect 38384 20674 38436 20680
rect 38396 20505 38424 20674
rect 38382 20496 38438 20505
rect 38382 20431 38438 20440
rect 37188 18352 37240 18358
rect 37188 18294 37240 18300
rect 37556 18080 37608 18086
rect 37556 18022 37608 18028
rect 35900 8900 35952 8906
rect 35900 8842 35952 8848
rect 36820 8900 36872 8906
rect 36820 8842 36872 8848
rect 35912 8566 35940 8842
rect 35900 8560 35952 8566
rect 35900 8502 35952 8508
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34428 6724 34480 6730
rect 34428 6666 34480 6672
rect 33140 6452 33192 6458
rect 33140 6394 33192 6400
rect 32588 6180 32640 6186
rect 32588 6122 32640 6128
rect 32772 6180 32824 6186
rect 32772 6122 32824 6128
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 32036 5908 32088 5914
rect 32036 5850 32088 5856
rect 32220 5908 32272 5914
rect 32220 5850 32272 5856
rect 32128 5704 32180 5710
rect 32128 5646 32180 5652
rect 31944 5636 31996 5642
rect 31944 5578 31996 5584
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 30656 5092 30708 5098
rect 30656 5034 30708 5040
rect 30288 5024 30340 5030
rect 30288 4966 30340 4972
rect 30196 4820 30248 4826
rect 30196 4762 30248 4768
rect 30300 4622 30328 4966
rect 30668 4758 30696 5034
rect 30656 4752 30708 4758
rect 30656 4694 30708 4700
rect 30288 4616 30340 4622
rect 30288 4558 30340 4564
rect 31772 4554 31800 5170
rect 31760 4548 31812 4554
rect 31760 4490 31812 4496
rect 31956 4486 31984 5578
rect 32140 5370 32168 5646
rect 32128 5364 32180 5370
rect 32128 5306 32180 5312
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 31944 4480 31996 4486
rect 31944 4422 31996 4428
rect 27896 4140 27948 4146
rect 27896 4082 27948 4088
rect 30104 4140 30156 4146
rect 30104 4082 30156 4088
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 37568 3126 37596 18022
rect 38384 18012 38436 18018
rect 38384 17954 38436 17960
rect 38396 17785 38424 17954
rect 38382 17776 38438 17785
rect 38382 17711 38438 17720
rect 37832 15904 37884 15910
rect 37832 15846 37884 15852
rect 37844 15745 37872 15846
rect 37830 15736 37886 15745
rect 37830 15671 37886 15680
rect 37924 11076 37976 11082
rect 37924 11018 37976 11024
rect 37936 10985 37964 11018
rect 37922 10976 37978 10985
rect 37922 10911 37978 10920
rect 38292 8968 38344 8974
rect 38290 8936 38292 8945
rect 38344 8936 38346 8945
rect 38290 8871 38346 8880
rect 37556 3120 37608 3126
rect 37556 3062 37608 3068
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 25964 3052 26016 3058
rect 25964 2994 26016 3000
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 37188 2848 37240 2854
rect 37188 2790 37240 2796
rect 14660 2746 14780 2774
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 32 800 60 2314
rect 2056 1170 2084 2314
rect 3988 1170 4016 2314
rect 6564 1170 6592 2314
rect 8496 1306 8524 2382
rect 14660 2378 14688 2746
rect 14936 2446 14964 2790
rect 17420 2446 17448 2790
rect 19812 2446 19840 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 19800 2440 19852 2446
rect 19800 2382 19852 2388
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 19432 2372 19484 2378
rect 19432 2314 19484 2320
rect 1964 1142 2084 1170
rect 3896 1142 4016 1170
rect 6472 1142 6592 1170
rect 8404 1278 8524 1306
rect 1964 800 1992 1142
rect 3896 800 3924 1142
rect 6472 800 6500 1142
rect 8404 800 8432 1278
rect 10980 800 11008 2314
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 12912 800 12940 2246
rect 15028 1170 15056 2246
rect 14844 1142 15056 1170
rect 14844 800 14872 1142
rect 17420 800 17448 2246
rect 19444 1170 19472 2314
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19352 1142 19472 1170
rect 19352 800 19380 1142
rect 26436 800 26464 2246
rect 37200 1465 37228 2790
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 37186 1456 37242 1465
rect 37186 1391 37242 1400
rect 37476 1306 37504 2382
rect 37384 1278 37504 1306
rect 37384 800 37412 1278
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 14830 0 14886 800
rect 17406 0 17462 800
rect 19338 0 19394 800
rect 21914 0 21970 800
rect 23846 0 23902 800
rect 26422 0 26478 800
rect 28354 0 28410 800
rect 30286 0 30342 800
rect 32862 0 32918 800
rect 34794 0 34850 800
rect 37370 0 37426 800
rect 39302 0 39358 800
<< via2 >>
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 938 36760 994 36816
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 5170 38392 5226 38448
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 938 25200 994 25256
rect 1490 20576 1546 20632
rect 938 18400 994 18456
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4066 27240 4122 27296
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 2962 22636 3018 22672
rect 2962 22616 2964 22636
rect 2964 22616 3016 22636
rect 3016 22616 3018 22636
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 938 15700 994 15736
rect 938 15680 940 15700
rect 940 15680 992 15700
rect 992 15680 994 15700
rect 1490 13640 1546 13696
rect 938 11600 994 11656
rect 938 8900 994 8936
rect 938 8880 940 8900
rect 940 8880 992 8900
rect 992 8880 994 8900
rect 1490 6840 1546 6896
rect 938 4120 994 4176
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4894 23060 4896 23080
rect 4896 23060 4948 23080
rect 4948 23060 4950 23080
rect 4894 23024 4950 23060
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 8298 29144 8354 29200
rect 6550 23296 6606 23352
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 3238 9580 3294 9616
rect 3238 9560 3240 9580
rect 3240 9560 3292 9580
rect 3292 9560 3294 9580
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4158 9016 4214 9072
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 5722 21120 5778 21176
rect 5630 20868 5686 20904
rect 5630 20848 5632 20868
rect 5632 20848 5684 20868
rect 5684 20848 5686 20868
rect 5998 18808 6054 18864
rect 7746 23296 7802 23352
rect 8022 23024 8078 23080
rect 7930 19352 7986 19408
rect 20350 38936 20406 38992
rect 8574 20168 8630 20224
rect 8390 19796 8392 19816
rect 8392 19796 8444 19816
rect 8444 19796 8446 19816
rect 8390 19760 8446 19796
rect 9034 20304 9090 20360
rect 9862 24112 9918 24168
rect 9678 21548 9734 21584
rect 9678 21528 9680 21548
rect 9680 21528 9732 21548
rect 9732 21528 9734 21548
rect 10046 21256 10102 21312
rect 9586 20712 9642 20768
rect 9494 19896 9550 19952
rect 9034 17856 9090 17912
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10138 20440 10194 20496
rect 11702 37748 11704 37768
rect 11704 37748 11756 37768
rect 11756 37748 11758 37768
rect 11702 37712 11758 37748
rect 10322 21548 10378 21584
rect 10322 21528 10324 21548
rect 10324 21528 10376 21548
rect 10376 21528 10378 21548
rect 10598 21528 10654 21584
rect 9586 14340 9642 14376
rect 9586 14320 9588 14340
rect 9588 14320 9640 14340
rect 9640 14320 9642 14340
rect 9586 13640 9642 13696
rect 11334 22480 11390 22536
rect 12070 32836 12126 32872
rect 12070 32816 12072 32836
rect 12072 32816 12124 32836
rect 12124 32816 12126 32836
rect 11518 28736 11574 28792
rect 12254 28736 12310 28792
rect 12346 25336 12402 25392
rect 10874 17992 10930 18048
rect 10230 12960 10286 13016
rect 11242 19080 11298 19136
rect 11334 15544 11390 15600
rect 15566 38664 15622 38720
rect 12530 37868 12586 37904
rect 12530 37848 12532 37868
rect 12532 37848 12584 37868
rect 12584 37848 12586 37868
rect 22374 38664 22430 38720
rect 27066 38664 27122 38720
rect 25778 38392 25834 38448
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 12990 31864 13046 31920
rect 12898 29028 12954 29064
rect 12898 29008 12900 29028
rect 12900 29008 12952 29028
rect 12952 29008 12954 29028
rect 13634 32000 13690 32056
rect 12622 23432 12678 23488
rect 11518 15408 11574 15464
rect 12898 19624 12954 19680
rect 12346 16108 12402 16144
rect 12346 16088 12348 16108
rect 12348 16088 12400 16108
rect 12400 16088 12402 16108
rect 12254 15952 12310 16008
rect 12162 8472 12218 8528
rect 14278 33768 14334 33824
rect 14738 33904 14794 33960
rect 13910 28872 13966 28928
rect 14830 27920 14886 27976
rect 13726 24384 13782 24440
rect 13726 23604 13728 23624
rect 13728 23604 13780 23624
rect 13780 23604 13782 23624
rect 13726 23568 13782 23604
rect 13726 21392 13782 21448
rect 13726 19488 13782 19544
rect 14186 25880 14242 25936
rect 14738 26988 14794 27024
rect 14738 26968 14740 26988
rect 14740 26968 14792 26988
rect 14792 26968 14794 26988
rect 14278 23740 14280 23760
rect 14280 23740 14332 23760
rect 14332 23740 14334 23760
rect 14278 23704 14334 23740
rect 15382 34060 15438 34096
rect 15382 34040 15384 34060
rect 15384 34040 15436 34060
rect 15436 34040 15438 34060
rect 15566 34312 15622 34368
rect 16486 34196 16542 34232
rect 16486 34176 16488 34196
rect 16488 34176 16540 34196
rect 16540 34176 16542 34196
rect 15842 31456 15898 31512
rect 15658 29688 15714 29744
rect 15106 29280 15162 29336
rect 15198 24792 15254 24848
rect 14186 20984 14242 21040
rect 14738 21684 14794 21720
rect 14738 21664 14740 21684
rect 14740 21664 14792 21684
rect 14792 21664 14794 21684
rect 14646 19488 14702 19544
rect 14738 18264 14794 18320
rect 14370 14476 14426 14512
rect 14370 14456 14372 14476
rect 14372 14456 14424 14476
rect 14424 14456 14426 14476
rect 15198 21664 15254 21720
rect 16302 31184 16358 31240
rect 16394 30232 16450 30288
rect 15934 26424 15990 26480
rect 16854 31320 16910 31376
rect 17406 35980 17408 36000
rect 17408 35980 17460 36000
rect 17460 35980 17462 36000
rect 17406 35944 17462 35980
rect 19154 37712 19210 37768
rect 16854 27512 16910 27568
rect 16486 27240 16542 27296
rect 16486 26288 16542 26344
rect 17682 33088 17738 33144
rect 17958 34448 18014 34504
rect 17958 34040 18014 34096
rect 17958 31884 18014 31920
rect 17958 31864 17960 31884
rect 17960 31864 18012 31884
rect 18012 31864 18014 31884
rect 17866 31456 17922 31512
rect 18418 32000 18474 32056
rect 17682 29688 17738 29744
rect 17682 28872 17738 28928
rect 15658 18672 15714 18728
rect 12530 3984 12586 4040
rect 13174 3984 13230 4040
rect 14922 8472 14978 8528
rect 16118 21664 16174 21720
rect 17314 26188 17316 26208
rect 17316 26188 17368 26208
rect 17368 26188 17370 26208
rect 17314 26152 17370 26188
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 18602 33924 18658 33960
rect 18602 33904 18604 33924
rect 18604 33904 18656 33924
rect 18656 33904 18658 33924
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 20166 35944 20222 36000
rect 20442 35944 20498 36000
rect 19890 35672 19946 35728
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19246 34176 19302 34232
rect 19154 34040 19210 34096
rect 19062 33224 19118 33280
rect 18694 32136 18750 32192
rect 18326 30368 18382 30424
rect 17958 29552 18014 29608
rect 18050 28872 18106 28928
rect 18050 28736 18106 28792
rect 17866 27532 17922 27568
rect 17866 27512 17868 27532
rect 17868 27512 17920 27532
rect 17920 27512 17922 27532
rect 17682 27240 17738 27296
rect 17682 26424 17738 26480
rect 17774 26152 17830 26208
rect 19338 33768 19394 33824
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19062 30776 19118 30832
rect 19246 30640 19302 30696
rect 18878 29008 18934 29064
rect 19154 29144 19210 29200
rect 17682 24248 17738 24304
rect 17314 23432 17370 23488
rect 17498 22516 17500 22536
rect 17500 22516 17552 22536
rect 17552 22516 17554 22536
rect 17498 22480 17554 22516
rect 17222 20032 17278 20088
rect 17222 19760 17278 19816
rect 18970 26988 19026 27024
rect 18970 26968 18972 26988
rect 18972 26968 19024 26988
rect 19024 26968 19026 26988
rect 18786 26288 18842 26344
rect 18694 25472 18750 25528
rect 18970 26424 19026 26480
rect 19154 28736 19210 28792
rect 20258 34312 20314 34368
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19522 29960 19578 30016
rect 19706 29824 19762 29880
rect 20074 30368 20130 30424
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19706 28872 19762 28928
rect 19522 28464 19578 28520
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19430 28056 19486 28112
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19154 24268 19210 24304
rect 19154 24248 19156 24268
rect 19156 24248 19208 24268
rect 19208 24248 19210 24268
rect 20258 30912 20314 30968
rect 21086 33496 21142 33552
rect 20626 33360 20682 33416
rect 20626 33224 20682 33280
rect 20718 31048 20774 31104
rect 21086 32816 21142 32872
rect 21730 33940 21732 33960
rect 21732 33940 21784 33960
rect 21784 33940 21786 33960
rect 21730 33904 21786 33940
rect 21270 32428 21326 32464
rect 21270 32408 21272 32428
rect 21272 32408 21324 32428
rect 21324 32408 21326 32428
rect 21270 31764 21272 31784
rect 21272 31764 21324 31784
rect 21324 31764 21326 31784
rect 21270 31728 21326 31764
rect 20350 30504 20406 30560
rect 20258 30096 20314 30152
rect 20166 29960 20222 30016
rect 20258 29416 20314 29472
rect 20534 30096 20590 30152
rect 20810 30232 20866 30288
rect 20258 28600 20314 28656
rect 20074 26288 20130 26344
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 20810 29280 20866 29336
rect 20994 29280 21050 29336
rect 20718 28192 20774 28248
rect 20258 25744 20314 25800
rect 20258 25336 20314 25392
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 18602 23432 18658 23488
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19522 23724 19578 23760
rect 19522 23704 19524 23724
rect 19524 23704 19576 23724
rect 19576 23704 19578 23724
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 21822 33516 21878 33552
rect 21822 33496 21824 33516
rect 21824 33496 21876 33516
rect 21876 33496 21878 33516
rect 22098 33260 22100 33280
rect 22100 33260 22152 33280
rect 22152 33260 22154 33280
rect 22098 33224 22154 33260
rect 21822 31456 21878 31512
rect 21546 31204 21602 31240
rect 21546 31184 21548 31204
rect 21548 31184 21600 31204
rect 21600 31184 21602 31204
rect 21362 30912 21418 30968
rect 21546 29416 21602 29472
rect 20902 27920 20958 27976
rect 20810 26424 20866 26480
rect 21178 27784 21234 27840
rect 21454 28872 21510 28928
rect 21638 29164 21694 29200
rect 21638 29144 21640 29164
rect 21640 29144 21692 29164
rect 21692 29144 21694 29164
rect 22558 34176 22614 34232
rect 22466 33804 22468 33824
rect 22468 33804 22520 33824
rect 22520 33804 22522 33824
rect 22466 33768 22522 33804
rect 22926 37324 22982 37360
rect 22926 37304 22928 37324
rect 22928 37304 22980 37324
rect 22980 37304 22982 37324
rect 22098 29008 22154 29064
rect 21454 25744 21510 25800
rect 21914 27648 21970 27704
rect 21822 26424 21878 26480
rect 23018 34040 23074 34096
rect 22926 33904 22982 33960
rect 22834 32852 22836 32872
rect 22836 32852 22888 32872
rect 22888 32852 22890 32872
rect 22834 32816 22890 32852
rect 22558 31864 22614 31920
rect 22742 31320 22798 31376
rect 23110 33904 23166 33960
rect 23202 33768 23258 33824
rect 23018 31340 23074 31376
rect 23018 31320 23020 31340
rect 23020 31320 23072 31340
rect 23072 31320 23074 31340
rect 22834 30368 22890 30424
rect 22742 29588 22744 29608
rect 22744 29588 22796 29608
rect 22796 29588 22798 29608
rect 22742 29552 22798 29588
rect 22558 28600 22614 28656
rect 21730 23704 21786 23760
rect 22098 24112 22154 24168
rect 18142 20576 18198 20632
rect 18050 18708 18052 18728
rect 18052 18708 18104 18728
rect 18104 18708 18106 18728
rect 18050 18672 18106 18708
rect 18234 18128 18290 18184
rect 18234 17856 18290 17912
rect 18418 18708 18420 18728
rect 18420 18708 18472 18728
rect 18472 18708 18474 18728
rect 18418 18672 18474 18708
rect 18418 17856 18474 17912
rect 17590 15544 17646 15600
rect 17774 14492 17776 14512
rect 17776 14492 17828 14512
rect 17828 14492 17830 14512
rect 17774 14456 17830 14492
rect 19062 20576 19118 20632
rect 19062 18300 19064 18320
rect 19064 18300 19116 18320
rect 19116 18300 19118 18320
rect 19062 18264 19118 18300
rect 18970 18128 19026 18184
rect 17498 10532 17554 10568
rect 17498 10512 17500 10532
rect 17500 10512 17552 10532
rect 17552 10512 17554 10532
rect 18694 12960 18750 13016
rect 18694 11620 18750 11656
rect 18694 11600 18696 11620
rect 18696 11600 18748 11620
rect 18748 11600 18750 11620
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 20074 21800 20130 21856
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19338 16496 19394 16552
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 18234 10376 18290 10432
rect 20350 20748 20352 20768
rect 20352 20748 20404 20768
rect 20404 20748 20406 20768
rect 20350 20712 20406 20748
rect 20994 21256 21050 21312
rect 21822 20712 21878 20768
rect 21914 20440 21970 20496
rect 22466 21836 22468 21856
rect 22468 21836 22520 21856
rect 22520 21836 22522 21856
rect 22466 21800 22522 21836
rect 22374 20884 22376 20904
rect 22376 20884 22428 20904
rect 22428 20884 22430 20904
rect 22374 20848 22430 20884
rect 22374 20304 22430 20360
rect 22098 19896 22154 19952
rect 22098 19216 22154 19272
rect 21454 17992 21510 18048
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 22374 19488 22430 19544
rect 22374 18944 22430 19000
rect 20810 10376 20866 10432
rect 23110 30504 23166 30560
rect 25318 37868 25374 37904
rect 25318 37848 25320 37868
rect 25320 37848 25372 37868
rect 25372 37848 25374 37868
rect 23478 34448 23534 34504
rect 23846 34604 23902 34640
rect 23846 34584 23848 34604
rect 23848 34584 23900 34604
rect 23900 34584 23902 34604
rect 23478 33396 23480 33416
rect 23480 33396 23532 33416
rect 23532 33396 23534 33416
rect 23478 33360 23534 33396
rect 23386 31456 23442 31512
rect 23386 29960 23442 30016
rect 24030 34176 24086 34232
rect 24030 33260 24032 33280
rect 24032 33260 24084 33280
rect 24084 33260 24086 33280
rect 24030 33224 24086 33260
rect 24306 33088 24362 33144
rect 23754 31048 23810 31104
rect 24306 31864 24362 31920
rect 25226 37304 25282 37360
rect 24030 31592 24086 31648
rect 23386 28736 23442 28792
rect 23570 29008 23626 29064
rect 23110 25900 23166 25936
rect 23110 25880 23112 25900
rect 23112 25880 23164 25900
rect 23164 25880 23166 25900
rect 22650 21664 22706 21720
rect 22650 17856 22706 17912
rect 22834 21392 22890 21448
rect 22926 21256 22982 21312
rect 23478 25472 23534 25528
rect 24214 28872 24270 28928
rect 24398 27784 24454 27840
rect 24306 25608 24362 25664
rect 23938 24384 23994 24440
rect 24306 23588 24362 23624
rect 24306 23568 24308 23588
rect 24308 23568 24360 23588
rect 24360 23568 24362 23588
rect 25134 30504 25190 30560
rect 24950 29824 25006 29880
rect 25134 26036 25190 26072
rect 25134 26016 25136 26036
rect 25136 26016 25188 26036
rect 25188 26016 25190 26036
rect 24950 25764 25006 25800
rect 24950 25744 24952 25764
rect 24952 25744 25004 25764
rect 25004 25744 25006 25764
rect 24858 22616 24914 22672
rect 24674 22072 24730 22128
rect 24858 21664 24914 21720
rect 23386 20168 23442 20224
rect 23478 19760 23534 19816
rect 23386 19624 23442 19680
rect 24858 21120 24914 21176
rect 25134 25472 25190 25528
rect 25042 21140 25098 21176
rect 25042 21120 25044 21140
rect 25044 21120 25096 21140
rect 25096 21120 25098 21140
rect 24030 19760 24086 19816
rect 23570 18808 23626 18864
rect 23386 17856 23442 17912
rect 23202 17584 23258 17640
rect 23294 16516 23350 16552
rect 23294 16496 23296 16516
rect 23296 16496 23348 16516
rect 23348 16496 23350 16516
rect 23754 15952 23810 16008
rect 24306 19252 24308 19272
rect 24308 19252 24360 19272
rect 24360 19252 24362 19272
rect 24306 19216 24362 19252
rect 23202 15020 23258 15056
rect 23202 15000 23204 15020
rect 23204 15000 23256 15020
rect 23256 15000 23258 15020
rect 21454 10956 21456 10976
rect 21456 10956 21508 10976
rect 21508 10956 21510 10976
rect 21454 10920 21510 10956
rect 21546 10648 21602 10704
rect 20350 9832 20406 9888
rect 18970 8492 19026 8528
rect 18970 8472 18972 8492
rect 18972 8472 19024 8492
rect 19024 8472 19026 8492
rect 18234 6840 18290 6896
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 22558 10920 22614 10976
rect 22282 9560 22338 9616
rect 23018 10648 23074 10704
rect 22834 9016 22890 9072
rect 23754 9288 23810 9344
rect 24950 19080 25006 19136
rect 25410 33260 25412 33280
rect 25412 33260 25464 33280
rect 25464 33260 25466 33280
rect 25410 33224 25466 33260
rect 25502 31728 25558 31784
rect 25410 26832 25466 26888
rect 25318 23160 25374 23216
rect 26790 33496 26846 33552
rect 26606 32000 26662 32056
rect 26606 31864 26662 31920
rect 26238 30504 26294 30560
rect 25962 29688 26018 29744
rect 26698 30368 26754 30424
rect 26238 28192 26294 28248
rect 26330 26968 26386 27024
rect 25870 26288 25926 26344
rect 26422 26424 26478 26480
rect 26330 25608 26386 25664
rect 25870 23704 25926 23760
rect 25962 23044 26018 23080
rect 25962 23024 25964 23044
rect 25964 23024 26016 23044
rect 26016 23024 26018 23044
rect 25870 21664 25926 21720
rect 25318 20576 25374 20632
rect 25318 19352 25374 19408
rect 25778 19488 25834 19544
rect 24674 17040 24730 17096
rect 24490 16496 24546 16552
rect 24490 16088 24546 16144
rect 24122 9832 24178 9888
rect 24490 9832 24546 9888
rect 23938 9152 23994 9208
rect 25134 15408 25190 15464
rect 24766 9288 24822 9344
rect 25502 9152 25558 9208
rect 21822 4564 21824 4584
rect 21824 4564 21876 4584
rect 21876 4564 21878 4584
rect 21822 4528 21878 4564
rect 25134 4528 25190 4584
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 25594 4564 25596 4584
rect 25596 4564 25648 4584
rect 25648 4564 25650 4584
rect 25594 4528 25650 4564
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 26054 21256 26110 21312
rect 26054 20032 26110 20088
rect 27986 37304 28042 37360
rect 27158 24792 27214 24848
rect 28446 35944 28502 36000
rect 28170 34448 28226 34504
rect 28446 34584 28502 34640
rect 27710 31084 27712 31104
rect 27712 31084 27764 31104
rect 27764 31084 27766 31104
rect 27710 31048 27766 31084
rect 27894 25472 27950 25528
rect 27710 23296 27766 23352
rect 27710 22072 27766 22128
rect 26330 19760 26386 19816
rect 26330 14864 26386 14920
rect 27710 21392 27766 21448
rect 27710 21120 27766 21176
rect 27894 21564 27896 21584
rect 27896 21564 27948 21584
rect 27948 21564 27950 21584
rect 27894 21528 27950 21564
rect 27342 19896 27398 19952
rect 27066 19388 27068 19408
rect 27068 19388 27120 19408
rect 27120 19388 27122 19408
rect 27066 19352 27122 19388
rect 27618 19488 27674 19544
rect 29274 31592 29330 31648
rect 28262 26832 28318 26888
rect 27894 19352 27950 19408
rect 27710 17740 27766 17776
rect 27710 17720 27712 17740
rect 27712 17720 27764 17740
rect 27764 17720 27766 17740
rect 28262 19372 28318 19408
rect 28262 19352 28264 19372
rect 28264 19352 28316 19372
rect 28316 19352 28318 19372
rect 28998 19896 29054 19952
rect 29274 26016 29330 26072
rect 29458 33088 29514 33144
rect 29090 19624 29146 19680
rect 26330 8780 26332 8800
rect 26332 8780 26384 8800
rect 26384 8780 26386 8800
rect 26330 8744 26386 8780
rect 27618 15156 27674 15192
rect 27618 15136 27620 15156
rect 27620 15136 27672 15156
rect 27672 15136 27674 15156
rect 27618 13368 27674 13424
rect 27710 11600 27766 11656
rect 27894 10512 27950 10568
rect 27986 10376 28042 10432
rect 26882 8880 26938 8936
rect 27802 8744 27858 8800
rect 27986 8916 27988 8936
rect 27988 8916 28040 8936
rect 28040 8916 28042 8936
rect 27986 8880 28042 8916
rect 28446 15136 28502 15192
rect 28722 15020 28778 15056
rect 28722 15000 28724 15020
rect 28724 15000 28776 15020
rect 28776 15000 28778 15020
rect 28538 14884 28594 14920
rect 28538 14864 28540 14884
rect 28540 14864 28592 14884
rect 28592 14864 28594 14884
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 37646 38820 37702 38856
rect 37646 38800 37648 38820
rect 37648 38800 37700 38820
rect 37700 38800 37702 38820
rect 37922 38800 37978 38856
rect 30194 30776 30250 30832
rect 29826 29688 29882 29744
rect 29918 27920 29974 27976
rect 30654 30796 30710 30832
rect 30654 30776 30656 30796
rect 30656 30776 30708 30796
rect 30708 30776 30710 30796
rect 30930 30660 30986 30696
rect 30930 30640 30932 30660
rect 30932 30640 30984 30660
rect 30984 30640 30986 30660
rect 30562 29280 30618 29336
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37830 36760 37886 36816
rect 31574 29552 31630 29608
rect 30470 26324 30472 26344
rect 30472 26324 30524 26344
rect 30524 26324 30526 26344
rect 30470 26288 30526 26324
rect 31574 26036 31630 26072
rect 31574 26016 31576 26036
rect 31576 26016 31628 26036
rect 31628 26016 31630 26036
rect 31390 25916 31392 25936
rect 31392 25916 31444 25936
rect 31444 25916 31446 25936
rect 31390 25880 31446 25916
rect 32494 26036 32550 26072
rect 32494 26016 32496 26036
rect 32496 26016 32548 26036
rect 32548 26016 32550 26036
rect 30654 19896 30710 19952
rect 30378 18300 30380 18320
rect 30380 18300 30432 18320
rect 30432 18300 30434 18320
rect 30378 18264 30434 18300
rect 31114 19352 31170 19408
rect 29182 16088 29238 16144
rect 29642 16124 29644 16144
rect 29644 16124 29696 16144
rect 29696 16124 29698 16144
rect 29642 16088 29698 16124
rect 28630 10376 28686 10432
rect 30194 14320 30250 14376
rect 30194 10104 30250 10160
rect 30010 9424 30066 9480
rect 30654 9424 30710 9480
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 32494 23160 32550 23216
rect 33782 32408 33838 32464
rect 33690 29552 33746 29608
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 37922 34040 37978 34096
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34058 30776 34114 30832
rect 33322 25900 33378 25936
rect 33322 25880 33324 25900
rect 33324 25880 33376 25900
rect 33376 25880 33378 25900
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 36266 29688 36322 29744
rect 36634 29688 36690 29744
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 32034 17176 32090 17232
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34610 21664 34666 21720
rect 33782 18264 33838 18320
rect 32862 17196 32918 17232
rect 32862 17176 32864 17196
rect 32864 17176 32916 17196
rect 32916 17176 32918 17196
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 37830 22500 37886 22536
rect 37830 22480 37832 22500
rect 37832 22480 37884 22500
rect 37884 22480 37886 22500
rect 36818 21392 36874 21448
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 32862 10104 32918 10160
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 38382 20440 38438 20496
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38382 17720 38438 17776
rect 37830 15680 37886 15736
rect 37922 10920 37978 10976
rect 38290 8916 38292 8936
rect 38292 8916 38344 8936
rect 38344 8916 38346 8936
rect 38290 8880 38346 8916
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 37186 1400 37242 1456
<< metal3 >>
rect 0 39448 800 39568
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 14222 38932 14228 38996
rect 14292 38994 14298 38996
rect 20345 38994 20411 38997
rect 14292 38992 20411 38994
rect 14292 38936 20350 38992
rect 20406 38936 20411 38992
rect 14292 38934 20411 38936
rect 14292 38932 14298 38934
rect 20345 38931 20411 38934
rect 9806 38796 9812 38860
rect 9876 38858 9882 38860
rect 37641 38858 37707 38861
rect 9876 38856 37707 38858
rect 9876 38800 37646 38856
rect 37702 38800 37707 38856
rect 9876 38798 37707 38800
rect 9876 38796 9882 38798
rect 37641 38795 37707 38798
rect 37917 38858 37983 38861
rect 38618 38858 39418 38888
rect 37917 38856 39418 38858
rect 37917 38800 37922 38856
rect 37978 38800 39418 38856
rect 37917 38798 39418 38800
rect 37917 38795 37983 38798
rect 38618 38768 39418 38798
rect 10358 38660 10364 38724
rect 10428 38722 10434 38724
rect 15561 38722 15627 38725
rect 10428 38720 15627 38722
rect 10428 38664 15566 38720
rect 15622 38664 15627 38720
rect 10428 38662 15627 38664
rect 10428 38660 10434 38662
rect 15561 38659 15627 38662
rect 22369 38722 22435 38725
rect 22870 38722 22876 38724
rect 22369 38720 22876 38722
rect 22369 38664 22374 38720
rect 22430 38664 22876 38720
rect 22369 38662 22876 38664
rect 22369 38659 22435 38662
rect 22870 38660 22876 38662
rect 22940 38660 22946 38724
rect 23974 38660 23980 38724
rect 24044 38722 24050 38724
rect 27061 38722 27127 38725
rect 24044 38720 27127 38722
rect 24044 38664 27066 38720
rect 27122 38664 27127 38720
rect 24044 38662 27127 38664
rect 24044 38660 24050 38662
rect 27061 38659 27127 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 5165 38450 5231 38453
rect 25773 38450 25839 38453
rect 5165 38448 25839 38450
rect 5165 38392 5170 38448
rect 5226 38392 25778 38448
rect 25834 38392 25839 38448
rect 5165 38390 25839 38392
rect 5165 38387 5231 38390
rect 25773 38387 25839 38390
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 12525 37906 12591 37909
rect 25313 37906 25379 37909
rect 12525 37904 25379 37906
rect 12525 37848 12530 37904
rect 12586 37848 25318 37904
rect 25374 37848 25379 37904
rect 12525 37846 25379 37848
rect 12525 37843 12591 37846
rect 25313 37843 25379 37846
rect 11697 37770 11763 37773
rect 19149 37770 19215 37773
rect 11697 37768 19215 37770
rect 11697 37712 11702 37768
rect 11758 37712 19154 37768
rect 19210 37712 19215 37768
rect 11697 37710 19215 37712
rect 11697 37707 11763 37710
rect 19149 37707 19215 37710
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 22134 37300 22140 37364
rect 22204 37362 22210 37364
rect 22921 37362 22987 37365
rect 22204 37360 22987 37362
rect 22204 37304 22926 37360
rect 22982 37304 22987 37360
rect 22204 37302 22987 37304
rect 22204 37300 22210 37302
rect 22921 37299 22987 37302
rect 25221 37364 25287 37365
rect 25221 37360 25268 37364
rect 25332 37362 25338 37364
rect 25221 37304 25226 37360
rect 25221 37300 25268 37304
rect 25332 37302 25378 37362
rect 25332 37300 25338 37302
rect 27838 37300 27844 37364
rect 27908 37362 27914 37364
rect 27981 37362 28047 37365
rect 27908 37360 28047 37362
rect 27908 37304 27986 37360
rect 28042 37304 28047 37360
rect 27908 37302 28047 37304
rect 27908 37300 27914 37302
rect 25221 37299 25287 37300
rect 27981 37299 28047 37302
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 0 36818 800 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 800 36758
rect 933 36755 999 36758
rect 37825 36818 37891 36821
rect 38618 36818 39418 36848
rect 37825 36816 39418 36818
rect 37825 36760 37830 36816
rect 37886 36760 39418 36816
rect 37825 36758 39418 36760
rect 37825 36755 37891 36758
rect 38618 36728 39418 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 17401 36002 17467 36005
rect 17534 36002 17540 36004
rect 17401 36000 17540 36002
rect 17401 35944 17406 36000
rect 17462 35944 17540 36000
rect 17401 35942 17540 35944
rect 17401 35939 17467 35942
rect 17534 35940 17540 35942
rect 17604 35940 17610 36004
rect 20161 36002 20227 36005
rect 20437 36004 20503 36005
rect 20294 36002 20300 36004
rect 20161 36000 20300 36002
rect 20161 35944 20166 36000
rect 20222 35944 20300 36000
rect 20161 35942 20300 35944
rect 20161 35939 20227 35942
rect 20294 35940 20300 35942
rect 20364 35940 20370 36004
rect 20437 36000 20484 36004
rect 20548 36002 20554 36004
rect 28441 36002 28507 36005
rect 28942 36002 28948 36004
rect 20437 35944 20442 36000
rect 20437 35940 20484 35944
rect 20548 35942 20594 36002
rect 28441 36000 28948 36002
rect 28441 35944 28446 36000
rect 28502 35944 28948 36000
rect 28441 35942 28948 35944
rect 20548 35940 20554 35942
rect 20437 35939 20503 35940
rect 28441 35939 28507 35942
rect 28942 35940 28948 35942
rect 29012 35940 29018 36004
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 14774 35668 14780 35732
rect 14844 35730 14850 35732
rect 19885 35730 19951 35733
rect 14844 35728 19951 35730
rect 14844 35672 19890 35728
rect 19946 35672 19951 35728
rect 14844 35670 19951 35672
rect 14844 35668 14850 35670
rect 19885 35667 19951 35670
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 0 34688 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 23841 34642 23907 34645
rect 28441 34642 28507 34645
rect 23841 34640 28507 34642
rect 23841 34584 23846 34640
rect 23902 34584 28446 34640
rect 28502 34584 28507 34640
rect 23841 34582 28507 34584
rect 23841 34579 23907 34582
rect 28441 34579 28507 34582
rect 17953 34506 18019 34509
rect 23473 34506 23539 34509
rect 28165 34506 28231 34509
rect 17953 34504 28231 34506
rect 17953 34448 17958 34504
rect 18014 34448 23478 34504
rect 23534 34448 28170 34504
rect 28226 34448 28231 34504
rect 17953 34446 28231 34448
rect 17953 34443 18019 34446
rect 23473 34443 23539 34446
rect 28165 34443 28231 34446
rect 15561 34370 15627 34373
rect 20253 34370 20319 34373
rect 15561 34368 20319 34370
rect 15561 34312 15566 34368
rect 15622 34312 20258 34368
rect 20314 34312 20319 34368
rect 15561 34310 20319 34312
rect 15561 34307 15627 34310
rect 20253 34307 20319 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 16481 34234 16547 34237
rect 19241 34234 19307 34237
rect 16481 34232 19307 34234
rect 16481 34176 16486 34232
rect 16542 34176 19246 34232
rect 19302 34176 19307 34232
rect 16481 34174 19307 34176
rect 16481 34171 16547 34174
rect 19241 34171 19307 34174
rect 22553 34234 22619 34237
rect 24025 34234 24091 34237
rect 22553 34232 24091 34234
rect 22553 34176 22558 34232
rect 22614 34176 24030 34232
rect 24086 34176 24091 34232
rect 22553 34174 24091 34176
rect 22553 34171 22619 34174
rect 24025 34171 24091 34174
rect 15377 34098 15443 34101
rect 17953 34098 18019 34101
rect 15377 34096 18019 34098
rect 15377 34040 15382 34096
rect 15438 34040 17958 34096
rect 18014 34040 18019 34096
rect 15377 34038 18019 34040
rect 15377 34035 15443 34038
rect 17953 34035 18019 34038
rect 19149 34098 19215 34101
rect 23013 34098 23079 34101
rect 19149 34096 23079 34098
rect 19149 34040 19154 34096
rect 19210 34040 23018 34096
rect 23074 34040 23079 34096
rect 19149 34038 23079 34040
rect 19149 34035 19215 34038
rect 23013 34035 23079 34038
rect 37917 34098 37983 34101
rect 38618 34098 39418 34128
rect 37917 34096 39418 34098
rect 37917 34040 37922 34096
rect 37978 34040 39418 34096
rect 37917 34038 39418 34040
rect 37917 34035 37983 34038
rect 38618 34008 39418 34038
rect 14733 33962 14799 33965
rect 18597 33962 18663 33965
rect 14733 33960 18663 33962
rect 14733 33904 14738 33960
rect 14794 33904 18602 33960
rect 18658 33904 18663 33960
rect 14733 33902 18663 33904
rect 14733 33899 14799 33902
rect 18597 33899 18663 33902
rect 21725 33962 21791 33965
rect 22921 33962 22987 33965
rect 21725 33960 22987 33962
rect 21725 33904 21730 33960
rect 21786 33904 22926 33960
rect 22982 33904 22987 33960
rect 21725 33902 22987 33904
rect 21725 33899 21791 33902
rect 22921 33899 22987 33902
rect 23105 33962 23171 33965
rect 26182 33962 26188 33964
rect 23105 33960 26188 33962
rect 23105 33904 23110 33960
rect 23166 33904 26188 33960
rect 23105 33902 26188 33904
rect 23105 33899 23171 33902
rect 26182 33900 26188 33902
rect 26252 33900 26258 33964
rect 14273 33826 14339 33829
rect 19333 33826 19399 33829
rect 14273 33824 19399 33826
rect 14273 33768 14278 33824
rect 14334 33768 19338 33824
rect 19394 33768 19399 33824
rect 14273 33766 19399 33768
rect 14273 33763 14339 33766
rect 19333 33763 19399 33766
rect 22461 33826 22527 33829
rect 23197 33826 23263 33829
rect 22461 33824 23263 33826
rect 22461 33768 22466 33824
rect 22522 33768 23202 33824
rect 23258 33768 23263 33824
rect 22461 33766 23263 33768
rect 22461 33763 22527 33766
rect 23197 33763 23263 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 21081 33554 21147 33557
rect 21214 33554 21220 33556
rect 21081 33552 21220 33554
rect 21081 33496 21086 33552
rect 21142 33496 21220 33552
rect 21081 33494 21220 33496
rect 21081 33491 21147 33494
rect 21214 33492 21220 33494
rect 21284 33492 21290 33556
rect 21817 33554 21883 33557
rect 26785 33554 26851 33557
rect 21817 33552 26851 33554
rect 21817 33496 21822 33552
rect 21878 33496 26790 33552
rect 26846 33496 26851 33552
rect 21817 33494 26851 33496
rect 21817 33491 21883 33494
rect 26785 33491 26851 33494
rect 20621 33418 20687 33421
rect 23473 33418 23539 33421
rect 20621 33416 23539 33418
rect 20621 33360 20626 33416
rect 20682 33360 23478 33416
rect 23534 33360 23539 33416
rect 20621 33358 23539 33360
rect 20621 33355 20687 33358
rect 23473 33355 23539 33358
rect 19057 33284 19123 33285
rect 19006 33282 19012 33284
rect 18966 33222 19012 33282
rect 19076 33280 19123 33284
rect 19118 33224 19123 33280
rect 19006 33220 19012 33222
rect 19076 33220 19123 33224
rect 19057 33219 19123 33220
rect 20621 33282 20687 33285
rect 22093 33282 22159 33285
rect 20621 33280 22159 33282
rect 20621 33224 20626 33280
rect 20682 33224 22098 33280
rect 22154 33224 22159 33280
rect 20621 33222 22159 33224
rect 20621 33219 20687 33222
rect 22093 33219 22159 33222
rect 24025 33282 24091 33285
rect 25405 33284 25471 33285
rect 24526 33282 24532 33284
rect 24025 33280 24532 33282
rect 24025 33224 24030 33280
rect 24086 33224 24532 33280
rect 24025 33222 24532 33224
rect 24025 33219 24091 33222
rect 24526 33220 24532 33222
rect 24596 33220 24602 33284
rect 25405 33280 25452 33284
rect 25516 33282 25522 33284
rect 25405 33224 25410 33280
rect 25405 33220 25452 33224
rect 25516 33222 25562 33282
rect 25516 33220 25522 33222
rect 25405 33219 25471 33220
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 17677 33146 17743 33149
rect 24301 33146 24367 33149
rect 17677 33144 24367 33146
rect 17677 33088 17682 33144
rect 17738 33088 24306 33144
rect 24362 33088 24367 33144
rect 17677 33086 24367 33088
rect 17677 33083 17743 33086
rect 24301 33083 24367 33086
rect 28942 33084 28948 33148
rect 29012 33146 29018 33148
rect 29453 33146 29519 33149
rect 29012 33144 29519 33146
rect 29012 33088 29458 33144
rect 29514 33088 29519 33144
rect 29012 33086 29519 33088
rect 29012 33084 29018 33086
rect 29453 33083 29519 33086
rect 12065 32874 12131 32877
rect 21081 32874 21147 32877
rect 22829 32874 22895 32877
rect 12065 32872 22895 32874
rect 12065 32816 12070 32872
rect 12126 32816 21086 32872
rect 21142 32816 22834 32872
rect 22890 32816 22895 32872
rect 12065 32814 22895 32816
rect 12065 32811 12131 32814
rect 21081 32811 21147 32814
rect 22829 32811 22895 32814
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 21265 32466 21331 32469
rect 33777 32466 33843 32469
rect 21265 32464 33843 32466
rect 21265 32408 21270 32464
rect 21326 32408 33782 32464
rect 33838 32408 33843 32464
rect 21265 32406 33843 32408
rect 21265 32403 21331 32406
rect 33777 32403 33843 32406
rect 18086 32132 18092 32196
rect 18156 32194 18162 32196
rect 18689 32194 18755 32197
rect 18156 32192 18755 32194
rect 18156 32136 18694 32192
rect 18750 32136 18755 32192
rect 18156 32134 18755 32136
rect 18156 32132 18162 32134
rect 18689 32131 18755 32134
rect 4210 32128 4526 32129
rect 0 31968 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 13629 32058 13695 32061
rect 15694 32058 15700 32060
rect 13629 32056 15700 32058
rect 13629 32000 13634 32056
rect 13690 32000 15700 32056
rect 13629 31998 15700 32000
rect 13629 31995 13695 31998
rect 15694 31996 15700 31998
rect 15764 31996 15770 32060
rect 18270 31996 18276 32060
rect 18340 32058 18346 32060
rect 18413 32058 18479 32061
rect 26601 32058 26667 32061
rect 28942 32058 28948 32060
rect 18340 32056 18479 32058
rect 18340 32000 18418 32056
rect 18474 32000 18479 32056
rect 18340 31998 18479 32000
rect 18340 31996 18346 31998
rect 18413 31995 18479 31998
rect 22050 32056 28948 32058
rect 22050 32000 26606 32056
rect 26662 32000 28948 32056
rect 22050 31998 28948 32000
rect 12985 31922 13051 31925
rect 17953 31922 18019 31925
rect 22050 31922 22110 31998
rect 26601 31995 26667 31998
rect 28942 31996 28948 31998
rect 29012 31996 29018 32060
rect 38618 31968 39418 32088
rect 12985 31920 22110 31922
rect 12985 31864 12990 31920
rect 13046 31864 17958 31920
rect 18014 31864 22110 31920
rect 12985 31862 22110 31864
rect 22553 31922 22619 31925
rect 24301 31922 24367 31925
rect 26601 31922 26667 31925
rect 22553 31920 26667 31922
rect 22553 31864 22558 31920
rect 22614 31864 24306 31920
rect 24362 31864 26606 31920
rect 26662 31864 26667 31920
rect 22553 31862 26667 31864
rect 12985 31859 13051 31862
rect 17953 31859 18019 31862
rect 22553 31859 22619 31862
rect 24301 31859 24367 31862
rect 26601 31859 26667 31862
rect 21265 31786 21331 31789
rect 25497 31786 25563 31789
rect 21265 31784 25563 31786
rect 21265 31728 21270 31784
rect 21326 31728 25502 31784
rect 25558 31728 25563 31784
rect 21265 31726 25563 31728
rect 21265 31723 21331 31726
rect 25497 31723 25563 31726
rect 24025 31650 24091 31653
rect 29269 31650 29335 31653
rect 24025 31648 29335 31650
rect 24025 31592 24030 31648
rect 24086 31592 29274 31648
rect 29330 31592 29335 31648
rect 24025 31590 29335 31592
rect 24025 31587 24091 31590
rect 29269 31587 29335 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 15837 31514 15903 31517
rect 17861 31514 17927 31517
rect 15837 31512 17927 31514
rect 15837 31456 15842 31512
rect 15898 31456 17866 31512
rect 17922 31456 17927 31512
rect 15837 31454 17927 31456
rect 15837 31451 15903 31454
rect 17861 31451 17927 31454
rect 21817 31514 21883 31517
rect 23381 31514 23447 31517
rect 21817 31512 23447 31514
rect 21817 31456 21822 31512
rect 21878 31456 23386 31512
rect 23442 31456 23447 31512
rect 21817 31454 23447 31456
rect 21817 31451 21883 31454
rect 23381 31451 23447 31454
rect 16849 31378 16915 31381
rect 21214 31378 21220 31380
rect 16849 31376 21220 31378
rect 16849 31320 16854 31376
rect 16910 31320 21220 31376
rect 16849 31318 21220 31320
rect 16849 31315 16915 31318
rect 21214 31316 21220 31318
rect 21284 31316 21290 31380
rect 22737 31378 22803 31381
rect 23013 31378 23079 31381
rect 22737 31376 23079 31378
rect 22737 31320 22742 31376
rect 22798 31320 23018 31376
rect 23074 31320 23079 31376
rect 22737 31318 23079 31320
rect 22737 31315 22803 31318
rect 23013 31315 23079 31318
rect 16297 31242 16363 31245
rect 21541 31242 21607 31245
rect 16297 31240 21607 31242
rect 16297 31184 16302 31240
rect 16358 31184 21546 31240
rect 21602 31184 21607 31240
rect 16297 31182 21607 31184
rect 16297 31179 16363 31182
rect 21541 31179 21607 31182
rect 20713 31106 20779 31109
rect 23749 31106 23815 31109
rect 20713 31104 23815 31106
rect 20713 31048 20718 31104
rect 20774 31048 23754 31104
rect 23810 31048 23815 31104
rect 20713 31046 23815 31048
rect 20713 31043 20779 31046
rect 23749 31043 23815 31046
rect 27705 31106 27771 31109
rect 27838 31106 27844 31108
rect 27705 31104 27844 31106
rect 27705 31048 27710 31104
rect 27766 31048 27844 31104
rect 27705 31046 27844 31048
rect 27705 31043 27771 31046
rect 27838 31044 27844 31046
rect 27908 31044 27914 31108
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 20253 30970 20319 30973
rect 21357 30970 21423 30973
rect 20253 30968 21423 30970
rect 20253 30912 20258 30968
rect 20314 30912 21362 30968
rect 21418 30912 21423 30968
rect 20253 30910 21423 30912
rect 20253 30907 20319 30910
rect 21357 30907 21423 30910
rect 19057 30834 19123 30837
rect 30189 30834 30255 30837
rect 19057 30832 30255 30834
rect 19057 30776 19062 30832
rect 19118 30776 30194 30832
rect 30250 30776 30255 30832
rect 19057 30774 30255 30776
rect 19057 30771 19123 30774
rect 30189 30771 30255 30774
rect 30649 30834 30715 30837
rect 34053 30834 34119 30837
rect 30649 30832 34119 30834
rect 30649 30776 30654 30832
rect 30710 30776 34058 30832
rect 34114 30776 34119 30832
rect 30649 30774 34119 30776
rect 30649 30771 30715 30774
rect 34053 30771 34119 30774
rect 19241 30698 19307 30701
rect 30925 30698 30991 30701
rect 19241 30696 30991 30698
rect 19241 30640 19246 30696
rect 19302 30640 30930 30696
rect 30986 30640 30991 30696
rect 19241 30638 30991 30640
rect 19241 30635 19307 30638
rect 30925 30635 30991 30638
rect 20345 30562 20411 30565
rect 23105 30562 23171 30565
rect 20345 30560 23171 30562
rect 20345 30504 20350 30560
rect 20406 30504 23110 30560
rect 23166 30504 23171 30560
rect 20345 30502 23171 30504
rect 20345 30499 20411 30502
rect 23105 30499 23171 30502
rect 25129 30562 25195 30565
rect 26233 30562 26299 30565
rect 25129 30560 26299 30562
rect 25129 30504 25134 30560
rect 25190 30504 26238 30560
rect 26294 30504 26299 30560
rect 25129 30502 26299 30504
rect 25129 30499 25195 30502
rect 26233 30499 26299 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 18321 30426 18387 30429
rect 18454 30426 18460 30428
rect 18321 30424 18460 30426
rect 18321 30368 18326 30424
rect 18382 30368 18460 30424
rect 18321 30366 18460 30368
rect 18321 30363 18387 30366
rect 18454 30364 18460 30366
rect 18524 30364 18530 30428
rect 20069 30426 20135 30429
rect 20348 30426 20408 30499
rect 20069 30424 20408 30426
rect 20069 30368 20074 30424
rect 20130 30368 20408 30424
rect 20069 30366 20408 30368
rect 22829 30426 22895 30429
rect 26693 30428 26759 30429
rect 23974 30426 23980 30428
rect 22829 30424 23980 30426
rect 22829 30368 22834 30424
rect 22890 30368 23980 30424
rect 22829 30366 23980 30368
rect 20069 30363 20135 30366
rect 22829 30363 22895 30366
rect 23974 30364 23980 30366
rect 24044 30364 24050 30428
rect 26693 30424 26740 30428
rect 26804 30426 26810 30428
rect 26693 30368 26698 30424
rect 26693 30364 26740 30368
rect 26804 30366 26850 30426
rect 26804 30364 26810 30366
rect 26693 30363 26759 30364
rect 16389 30290 16455 30293
rect 20805 30290 20871 30293
rect 16389 30288 20871 30290
rect 16389 30232 16394 30288
rect 16450 30232 20810 30288
rect 20866 30232 20871 30288
rect 16389 30230 20871 30232
rect 16389 30227 16455 30230
rect 20805 30227 20871 30230
rect 20253 30154 20319 30157
rect 20529 30154 20595 30157
rect 20253 30152 20595 30154
rect 20253 30096 20258 30152
rect 20314 30096 20534 30152
rect 20590 30096 20595 30152
rect 20253 30094 20595 30096
rect 20253 30091 20319 30094
rect 20529 30091 20595 30094
rect 0 29928 800 30048
rect 19517 30018 19583 30021
rect 20161 30018 20227 30021
rect 23381 30018 23447 30021
rect 19517 30016 23447 30018
rect 19517 29960 19522 30016
rect 19578 29960 20166 30016
rect 20222 29960 23386 30016
rect 23442 29960 23447 30016
rect 19517 29958 23447 29960
rect 19517 29955 19583 29958
rect 20161 29955 20227 29958
rect 23381 29955 23447 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19701 29882 19767 29885
rect 24945 29882 25011 29885
rect 19701 29880 25011 29882
rect 19701 29824 19706 29880
rect 19762 29824 24950 29880
rect 25006 29824 25011 29880
rect 19701 29822 25011 29824
rect 19701 29819 19767 29822
rect 24945 29819 25011 29822
rect 15653 29746 15719 29749
rect 17677 29746 17743 29749
rect 25957 29746 26023 29749
rect 29821 29746 29887 29749
rect 36261 29746 36327 29749
rect 36629 29746 36695 29749
rect 15653 29744 29010 29746
rect 15653 29688 15658 29744
rect 15714 29688 17682 29744
rect 17738 29688 25962 29744
rect 26018 29688 29010 29744
rect 15653 29686 29010 29688
rect 15653 29683 15719 29686
rect 17677 29683 17743 29686
rect 25957 29683 26023 29686
rect 17953 29610 18019 29613
rect 22737 29610 22803 29613
rect 17953 29608 20178 29610
rect 17953 29552 17958 29608
rect 18014 29552 20178 29608
rect 17953 29550 20178 29552
rect 17953 29547 18019 29550
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 15101 29338 15167 29341
rect 20118 29338 20178 29550
rect 21038 29608 22803 29610
rect 21038 29552 22742 29608
rect 22798 29552 22803 29608
rect 21038 29550 22803 29552
rect 28950 29610 29010 29686
rect 29821 29744 36695 29746
rect 29821 29688 29826 29744
rect 29882 29688 36266 29744
rect 36322 29688 36634 29744
rect 36690 29688 36695 29744
rect 29821 29686 36695 29688
rect 29821 29683 29887 29686
rect 36261 29683 36327 29686
rect 36629 29683 36695 29686
rect 31569 29610 31635 29613
rect 33685 29610 33751 29613
rect 28950 29608 33751 29610
rect 28950 29552 31574 29608
rect 31630 29552 33690 29608
rect 33746 29552 33751 29608
rect 28950 29550 33751 29552
rect 20253 29474 20319 29477
rect 21038 29474 21098 29550
rect 22737 29547 22803 29550
rect 31569 29547 31635 29550
rect 33685 29547 33751 29550
rect 20253 29472 21098 29474
rect 20253 29416 20258 29472
rect 20314 29416 21098 29472
rect 20253 29414 21098 29416
rect 20253 29411 20319 29414
rect 21214 29412 21220 29476
rect 21284 29474 21290 29476
rect 21541 29474 21607 29477
rect 21284 29472 21607 29474
rect 21284 29416 21546 29472
rect 21602 29416 21607 29472
rect 21284 29414 21607 29416
rect 21284 29412 21290 29414
rect 21541 29411 21607 29414
rect 20805 29338 20871 29341
rect 15101 29336 19442 29338
rect 15101 29280 15106 29336
rect 15162 29280 19442 29336
rect 15101 29278 19442 29280
rect 20118 29336 20871 29338
rect 20118 29280 20810 29336
rect 20866 29280 20871 29336
rect 20118 29278 20871 29280
rect 15101 29275 15167 29278
rect 8293 29202 8359 29205
rect 19149 29202 19215 29205
rect 8293 29200 19215 29202
rect 8293 29144 8298 29200
rect 8354 29144 19154 29200
rect 19210 29144 19215 29200
rect 8293 29142 19215 29144
rect 19382 29202 19442 29278
rect 20805 29275 20871 29278
rect 20989 29338 21055 29341
rect 30557 29338 30623 29341
rect 20989 29336 30623 29338
rect 20989 29280 20994 29336
rect 21050 29280 30562 29336
rect 30618 29280 30623 29336
rect 20989 29278 30623 29280
rect 20989 29275 21055 29278
rect 30557 29275 30623 29278
rect 38618 29248 39418 29368
rect 21633 29202 21699 29205
rect 19382 29200 21699 29202
rect 19382 29144 21638 29200
rect 21694 29144 21699 29200
rect 19382 29142 21699 29144
rect 8293 29139 8359 29142
rect 19149 29139 19215 29142
rect 21633 29139 21699 29142
rect 12893 29066 12959 29069
rect 13302 29066 13308 29068
rect 12893 29064 13308 29066
rect 12893 29008 12898 29064
rect 12954 29008 13308 29064
rect 12893 29006 13308 29008
rect 12893 29003 12959 29006
rect 13302 29004 13308 29006
rect 13372 29004 13378 29068
rect 16430 29004 16436 29068
rect 16500 29066 16506 29068
rect 18873 29066 18939 29069
rect 22093 29066 22159 29069
rect 16500 29064 18939 29066
rect 16500 29008 18878 29064
rect 18934 29008 18939 29064
rect 16500 29006 18939 29008
rect 16500 29004 16506 29006
rect 18873 29003 18939 29006
rect 19014 29064 22159 29066
rect 19014 29008 22098 29064
rect 22154 29008 22159 29064
rect 19014 29006 22159 29008
rect 13905 28930 13971 28933
rect 17677 28930 17743 28933
rect 13905 28928 17743 28930
rect 13905 28872 13910 28928
rect 13966 28872 17682 28928
rect 17738 28872 17743 28928
rect 13905 28870 17743 28872
rect 13905 28867 13971 28870
rect 17677 28867 17743 28870
rect 18045 28930 18111 28933
rect 19014 28930 19074 29006
rect 22093 29003 22159 29006
rect 23565 29068 23631 29069
rect 23565 29064 23612 29068
rect 23676 29066 23682 29068
rect 23565 29008 23570 29064
rect 23565 29004 23612 29008
rect 23676 29006 23722 29066
rect 23676 29004 23682 29006
rect 23565 29003 23631 29004
rect 18045 28928 19074 28930
rect 18045 28872 18050 28928
rect 18106 28872 19074 28928
rect 18045 28870 19074 28872
rect 19701 28930 19767 28933
rect 21449 28930 21515 28933
rect 24209 28930 24275 28933
rect 19701 28928 24275 28930
rect 19701 28872 19706 28928
rect 19762 28872 21454 28928
rect 21510 28872 24214 28928
rect 24270 28872 24275 28928
rect 19701 28870 24275 28872
rect 18045 28867 18111 28870
rect 19701 28867 19767 28870
rect 21449 28867 21515 28870
rect 24209 28867 24275 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 11513 28794 11579 28797
rect 12249 28794 12315 28797
rect 18045 28796 18111 28797
rect 18045 28794 18092 28796
rect 11513 28792 18092 28794
rect 11513 28736 11518 28792
rect 11574 28736 12254 28792
rect 12310 28736 18050 28792
rect 11513 28734 18092 28736
rect 11513 28731 11579 28734
rect 12249 28731 12315 28734
rect 18045 28732 18092 28734
rect 18156 28732 18162 28796
rect 19149 28794 19215 28797
rect 23381 28794 23447 28797
rect 19149 28792 23447 28794
rect 19149 28736 19154 28792
rect 19210 28736 23386 28792
rect 23442 28736 23447 28792
rect 19149 28734 23447 28736
rect 18045 28731 18111 28732
rect 19149 28731 19215 28734
rect 23381 28731 23447 28734
rect 20253 28660 20319 28661
rect 20253 28658 20300 28660
rect 20172 28656 20300 28658
rect 20364 28658 20370 28660
rect 22553 28658 22619 28661
rect 20364 28656 22619 28658
rect 20172 28600 20258 28656
rect 20364 28600 22558 28656
rect 22614 28600 22619 28656
rect 20172 28598 20300 28600
rect 20253 28596 20300 28598
rect 20364 28598 22619 28600
rect 20364 28596 20370 28598
rect 20253 28595 20319 28596
rect 22553 28595 22619 28598
rect 19517 28522 19583 28525
rect 19382 28520 19583 28522
rect 19382 28464 19522 28520
rect 19578 28464 19583 28520
rect 19382 28462 19583 28464
rect 19382 28117 19442 28462
rect 19517 28459 19583 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 20713 28250 20779 28253
rect 25814 28250 25820 28252
rect 20713 28248 25820 28250
rect 20713 28192 20718 28248
rect 20774 28192 25820 28248
rect 20713 28190 25820 28192
rect 20713 28187 20779 28190
rect 25814 28188 25820 28190
rect 25884 28250 25890 28252
rect 26233 28250 26299 28253
rect 25884 28248 26299 28250
rect 25884 28192 26238 28248
rect 26294 28192 26299 28248
rect 25884 28190 26299 28192
rect 25884 28188 25890 28190
rect 26233 28187 26299 28190
rect 19382 28112 19491 28117
rect 19382 28056 19430 28112
rect 19486 28056 19491 28112
rect 19382 28054 19491 28056
rect 19425 28051 19491 28054
rect 14825 27978 14891 27981
rect 20897 27978 20963 27981
rect 14825 27976 20963 27978
rect 14825 27920 14830 27976
rect 14886 27920 20902 27976
rect 20958 27920 20963 27976
rect 14825 27918 20963 27920
rect 14825 27915 14891 27918
rect 20897 27915 20963 27918
rect 28942 27916 28948 27980
rect 29012 27978 29018 27980
rect 29913 27978 29979 27981
rect 29012 27976 29979 27978
rect 29012 27920 29918 27976
rect 29974 27920 29979 27976
rect 29012 27918 29979 27920
rect 29012 27916 29018 27918
rect 29913 27915 29979 27918
rect 21173 27842 21239 27845
rect 24393 27842 24459 27845
rect 21173 27840 24459 27842
rect 21173 27784 21178 27840
rect 21234 27784 24398 27840
rect 24454 27784 24459 27840
rect 21173 27782 24459 27784
rect 21173 27779 21239 27782
rect 24393 27779 24459 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 21909 27708 21975 27709
rect 21909 27704 21956 27708
rect 22020 27706 22026 27708
rect 21909 27648 21914 27704
rect 21909 27644 21956 27648
rect 22020 27646 22066 27706
rect 22020 27644 22026 27646
rect 21909 27643 21975 27644
rect 16849 27570 16915 27573
rect 17861 27570 17927 27573
rect 16849 27568 17927 27570
rect 16849 27512 16854 27568
rect 16910 27512 17866 27568
rect 17922 27512 17927 27568
rect 16849 27510 17927 27512
rect 16849 27507 16915 27510
rect 17861 27507 17927 27510
rect 0 27298 800 27328
rect 4061 27298 4127 27301
rect 0 27296 4127 27298
rect 0 27240 4066 27296
rect 4122 27240 4127 27296
rect 0 27238 4127 27240
rect 0 27208 800 27238
rect 4061 27235 4127 27238
rect 16481 27298 16547 27301
rect 17677 27298 17743 27301
rect 16481 27296 17743 27298
rect 16481 27240 16486 27296
rect 16542 27240 17682 27296
rect 17738 27240 17743 27296
rect 16481 27238 17743 27240
rect 16481 27235 16547 27238
rect 17677 27235 17743 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 38618 27208 39418 27328
rect 19570 27167 19886 27168
rect 14733 27026 14799 27029
rect 18965 27026 19031 27029
rect 26325 27026 26391 27029
rect 14733 27024 26391 27026
rect 14733 26968 14738 27024
rect 14794 26968 18970 27024
rect 19026 26968 26330 27024
rect 26386 26968 26391 27024
rect 14733 26966 26391 26968
rect 14733 26963 14799 26966
rect 18965 26963 19031 26966
rect 26325 26963 26391 26966
rect 25405 26890 25471 26893
rect 28257 26890 28323 26893
rect 25405 26888 28323 26890
rect 25405 26832 25410 26888
rect 25466 26832 28262 26888
rect 28318 26832 28323 26888
rect 25405 26830 28323 26832
rect 25405 26827 25471 26830
rect 28257 26827 28323 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 15929 26482 15995 26485
rect 17677 26482 17743 26485
rect 15929 26480 17743 26482
rect 15929 26424 15934 26480
rect 15990 26424 17682 26480
rect 17738 26424 17743 26480
rect 15929 26422 17743 26424
rect 15929 26419 15995 26422
rect 17677 26419 17743 26422
rect 18965 26482 19031 26485
rect 20805 26482 20871 26485
rect 18965 26480 20871 26482
rect 18965 26424 18970 26480
rect 19026 26424 20810 26480
rect 20866 26424 20871 26480
rect 18965 26422 20871 26424
rect 18965 26419 19031 26422
rect 20805 26419 20871 26422
rect 21817 26482 21883 26485
rect 26417 26482 26483 26485
rect 21817 26480 26483 26482
rect 21817 26424 21822 26480
rect 21878 26424 26422 26480
rect 26478 26424 26483 26480
rect 21817 26422 26483 26424
rect 21817 26419 21883 26422
rect 26417 26419 26483 26422
rect 16481 26346 16547 26349
rect 18781 26346 18847 26349
rect 16481 26344 18847 26346
rect 16481 26288 16486 26344
rect 16542 26288 18786 26344
rect 18842 26288 18847 26344
rect 16481 26286 18847 26288
rect 16481 26283 16547 26286
rect 18781 26283 18847 26286
rect 20069 26348 20135 26349
rect 20069 26344 20116 26348
rect 20180 26346 20186 26348
rect 25865 26346 25931 26349
rect 30465 26346 30531 26349
rect 20069 26288 20074 26344
rect 20069 26284 20116 26288
rect 20180 26286 20226 26346
rect 25865 26344 30531 26346
rect 25865 26288 25870 26344
rect 25926 26288 30470 26344
rect 30526 26288 30531 26344
rect 25865 26286 30531 26288
rect 20180 26284 20186 26286
rect 20069 26283 20135 26284
rect 25865 26283 25931 26286
rect 30465 26283 30531 26286
rect 17309 26210 17375 26213
rect 17769 26210 17835 26213
rect 17309 26208 17835 26210
rect 17309 26152 17314 26208
rect 17370 26152 17774 26208
rect 17830 26152 17835 26208
rect 17309 26150 17835 26152
rect 17309 26147 17375 26150
rect 17769 26147 17835 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 25129 26074 25195 26077
rect 25262 26074 25268 26076
rect 25129 26072 25268 26074
rect 25129 26016 25134 26072
rect 25190 26016 25268 26072
rect 25129 26014 25268 26016
rect 25129 26011 25195 26014
rect 25262 26012 25268 26014
rect 25332 26012 25338 26076
rect 29269 26074 29335 26077
rect 31569 26074 31635 26077
rect 32489 26074 32555 26077
rect 29269 26072 32555 26074
rect 29269 26016 29274 26072
rect 29330 26016 31574 26072
rect 31630 26016 32494 26072
rect 32550 26016 32555 26072
rect 29269 26014 32555 26016
rect 29269 26011 29335 26014
rect 31569 26011 31635 26014
rect 32489 26011 32555 26014
rect 14181 25938 14247 25941
rect 23105 25938 23171 25941
rect 14181 25936 23171 25938
rect 14181 25880 14186 25936
rect 14242 25880 23110 25936
rect 23166 25880 23171 25936
rect 14181 25878 23171 25880
rect 14181 25875 14247 25878
rect 23105 25875 23171 25878
rect 31385 25938 31451 25941
rect 33317 25938 33383 25941
rect 31385 25936 33383 25938
rect 31385 25880 31390 25936
rect 31446 25880 33322 25936
rect 33378 25880 33383 25936
rect 31385 25878 33383 25880
rect 31385 25875 31451 25878
rect 33317 25875 33383 25878
rect 20253 25802 20319 25805
rect 20478 25802 20484 25804
rect 20253 25800 20484 25802
rect 20253 25744 20258 25800
rect 20314 25744 20484 25800
rect 20253 25742 20484 25744
rect 20253 25739 20319 25742
rect 20478 25740 20484 25742
rect 20548 25740 20554 25804
rect 21449 25802 21515 25805
rect 24945 25802 25011 25805
rect 21449 25800 25011 25802
rect 21449 25744 21454 25800
rect 21510 25744 24950 25800
rect 25006 25744 25011 25800
rect 21449 25742 25011 25744
rect 21449 25739 21515 25742
rect 24945 25739 25011 25742
rect 24301 25666 24367 25669
rect 26325 25666 26391 25669
rect 24301 25664 26391 25666
rect 24301 25608 24306 25664
rect 24362 25608 26330 25664
rect 26386 25608 26391 25664
rect 24301 25606 26391 25608
rect 24301 25603 24367 25606
rect 26325 25603 26391 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 18689 25530 18755 25533
rect 23473 25530 23539 25533
rect 18689 25528 23539 25530
rect 18689 25472 18694 25528
rect 18750 25472 23478 25528
rect 23534 25472 23539 25528
rect 18689 25470 23539 25472
rect 18689 25467 18755 25470
rect 23473 25467 23539 25470
rect 25129 25530 25195 25533
rect 27889 25530 27955 25533
rect 25129 25528 27955 25530
rect 25129 25472 25134 25528
rect 25190 25472 27894 25528
rect 27950 25472 27955 25528
rect 25129 25470 27955 25472
rect 25129 25467 25195 25470
rect 27889 25467 27955 25470
rect 12341 25394 12407 25397
rect 20253 25394 20319 25397
rect 12341 25392 20319 25394
rect 12341 25336 12346 25392
rect 12402 25336 20258 25392
rect 20314 25336 20319 25392
rect 12341 25334 20319 25336
rect 12341 25331 12407 25334
rect 20253 25331 20319 25334
rect 0 25258 800 25288
rect 933 25258 999 25261
rect 0 25256 999 25258
rect 0 25200 938 25256
rect 994 25200 999 25256
rect 0 25198 999 25200
rect 0 25168 800 25198
rect 933 25195 999 25198
rect 38618 25168 39418 25288
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 15193 24850 15259 24853
rect 27153 24850 27219 24853
rect 15193 24848 27219 24850
rect 15193 24792 15198 24848
rect 15254 24792 27158 24848
rect 27214 24792 27219 24848
rect 15193 24790 27219 24792
rect 15193 24787 15259 24790
rect 27153 24787 27219 24790
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 13721 24442 13787 24445
rect 23933 24442 23999 24445
rect 13721 24440 23999 24442
rect 13721 24384 13726 24440
rect 13782 24384 23938 24440
rect 23994 24384 23999 24440
rect 13721 24382 23999 24384
rect 13721 24379 13787 24382
rect 23933 24379 23999 24382
rect 17677 24306 17743 24309
rect 19149 24306 19215 24309
rect 17677 24304 19215 24306
rect 17677 24248 17682 24304
rect 17738 24248 19154 24304
rect 19210 24248 19215 24304
rect 17677 24246 19215 24248
rect 17677 24243 17743 24246
rect 19149 24243 19215 24246
rect 9857 24170 9923 24173
rect 22093 24172 22159 24173
rect 22093 24170 22140 24172
rect 9857 24168 22140 24170
rect 22204 24170 22210 24172
rect 9857 24112 9862 24168
rect 9918 24112 22098 24168
rect 9857 24110 22140 24112
rect 9857 24107 9923 24110
rect 22093 24108 22140 24110
rect 22204 24110 22250 24170
rect 22204 24108 22210 24110
rect 22093 24107 22159 24108
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 14273 23762 14339 23765
rect 19517 23762 19583 23765
rect 21725 23762 21791 23765
rect 25865 23764 25931 23765
rect 14273 23760 21791 23762
rect 14273 23704 14278 23760
rect 14334 23704 19522 23760
rect 19578 23704 21730 23760
rect 21786 23704 21791 23760
rect 14273 23702 21791 23704
rect 14273 23699 14339 23702
rect 19517 23699 19583 23702
rect 21725 23699 21791 23702
rect 25814 23700 25820 23764
rect 25884 23762 25931 23764
rect 25884 23760 25976 23762
rect 25926 23704 25976 23760
rect 25884 23702 25976 23704
rect 25884 23700 25931 23702
rect 25865 23699 25931 23700
rect 13721 23626 13787 23629
rect 24301 23626 24367 23629
rect 13721 23624 24367 23626
rect 13721 23568 13726 23624
rect 13782 23568 24306 23624
rect 24362 23568 24367 23624
rect 13721 23566 24367 23568
rect 13721 23563 13787 23566
rect 24301 23563 24367 23566
rect 12617 23492 12683 23493
rect 12566 23490 12572 23492
rect 12526 23430 12572 23490
rect 12636 23488 12683 23492
rect 12678 23432 12683 23488
rect 12566 23428 12572 23430
rect 12636 23428 12683 23432
rect 12617 23427 12683 23428
rect 17309 23490 17375 23493
rect 18597 23490 18663 23493
rect 17309 23488 18663 23490
rect 17309 23432 17314 23488
rect 17370 23432 18602 23488
rect 18658 23432 18663 23488
rect 17309 23430 18663 23432
rect 17309 23427 17375 23430
rect 18597 23427 18663 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 6545 23354 6611 23357
rect 7741 23354 7807 23357
rect 27705 23354 27771 23357
rect 6545 23352 27771 23354
rect 6545 23296 6550 23352
rect 6606 23296 7746 23352
rect 7802 23296 27710 23352
rect 27766 23296 27771 23352
rect 6545 23294 27771 23296
rect 6545 23291 6611 23294
rect 7741 23291 7807 23294
rect 27705 23291 27771 23294
rect 0 23128 800 23248
rect 25313 23218 25379 23221
rect 32489 23218 32555 23221
rect 25313 23216 32555 23218
rect 25313 23160 25318 23216
rect 25374 23160 32494 23216
rect 32550 23160 32555 23216
rect 25313 23158 32555 23160
rect 25313 23155 25379 23158
rect 32489 23155 32555 23158
rect 4889 23082 4955 23085
rect 8017 23082 8083 23085
rect 25957 23082 26023 23085
rect 4889 23080 26023 23082
rect 4889 23024 4894 23080
rect 4950 23024 8022 23080
rect 8078 23024 25962 23080
rect 26018 23024 26023 23080
rect 4889 23022 26023 23024
rect 4889 23019 4955 23022
rect 8017 23019 8083 23022
rect 25957 23019 26023 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 2957 22674 3023 22677
rect 24853 22674 24919 22677
rect 2957 22672 24919 22674
rect 2957 22616 2962 22672
rect 3018 22616 24858 22672
rect 24914 22616 24919 22672
rect 2957 22614 24919 22616
rect 2957 22611 3023 22614
rect 24853 22611 24919 22614
rect 11329 22538 11395 22541
rect 17493 22538 17559 22541
rect 11329 22536 17559 22538
rect 11329 22480 11334 22536
rect 11390 22480 17498 22536
rect 17554 22480 17559 22536
rect 11329 22478 17559 22480
rect 11329 22475 11395 22478
rect 17493 22475 17559 22478
rect 37825 22538 37891 22541
rect 38618 22538 39418 22568
rect 37825 22536 39418 22538
rect 37825 22480 37830 22536
rect 37886 22480 39418 22536
rect 37825 22478 39418 22480
rect 37825 22475 37891 22478
rect 38618 22448 39418 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 24669 22130 24735 22133
rect 27705 22130 27771 22133
rect 24669 22128 27771 22130
rect 24669 22072 24674 22128
rect 24730 22072 27710 22128
rect 27766 22072 27771 22128
rect 24669 22070 27771 22072
rect 24669 22067 24735 22070
rect 27705 22067 27771 22070
rect 20069 21858 20135 21861
rect 22461 21858 22527 21861
rect 20069 21856 22527 21858
rect 20069 21800 20074 21856
rect 20130 21800 22466 21856
rect 22522 21800 22527 21856
rect 20069 21798 22527 21800
rect 20069 21795 20135 21798
rect 22461 21795 22527 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 14733 21724 14799 21725
rect 14733 21722 14780 21724
rect 14688 21720 14780 21722
rect 14688 21664 14738 21720
rect 14688 21662 14780 21664
rect 14733 21660 14780 21662
rect 14844 21660 14850 21724
rect 15193 21722 15259 21725
rect 16113 21722 16179 21725
rect 22645 21722 22711 21725
rect 15193 21720 16179 21722
rect 15193 21664 15198 21720
rect 15254 21664 16118 21720
rect 16174 21664 16179 21720
rect 15193 21662 16179 21664
rect 14733 21659 14799 21660
rect 15193 21659 15259 21662
rect 16113 21659 16179 21662
rect 22050 21720 22711 21722
rect 22050 21664 22650 21720
rect 22706 21664 22711 21720
rect 22050 21662 22711 21664
rect 9673 21586 9739 21589
rect 10317 21588 10383 21589
rect 9806 21586 9812 21588
rect 9673 21584 9812 21586
rect 9673 21528 9678 21584
rect 9734 21528 9812 21584
rect 9673 21526 9812 21528
rect 9673 21523 9739 21526
rect 9806 21524 9812 21526
rect 9876 21524 9882 21588
rect 10317 21586 10364 21588
rect 10272 21584 10364 21586
rect 10272 21528 10322 21584
rect 10272 21526 10364 21528
rect 10317 21524 10364 21526
rect 10428 21524 10434 21588
rect 10593 21586 10659 21589
rect 22050 21586 22110 21662
rect 22645 21659 22711 21662
rect 24853 21722 24919 21725
rect 25865 21722 25931 21725
rect 34605 21722 34671 21725
rect 24853 21720 34671 21722
rect 24853 21664 24858 21720
rect 24914 21664 25870 21720
rect 25926 21664 34610 21720
rect 34666 21664 34671 21720
rect 24853 21662 34671 21664
rect 24853 21659 24919 21662
rect 25865 21659 25931 21662
rect 34605 21659 34671 21662
rect 27889 21586 27955 21589
rect 10593 21584 22110 21586
rect 10593 21528 10598 21584
rect 10654 21528 22110 21584
rect 10593 21526 22110 21528
rect 22510 21584 27955 21586
rect 22510 21528 27894 21584
rect 27950 21528 27955 21584
rect 22510 21526 27955 21528
rect 10317 21523 10383 21524
rect 10593 21523 10659 21526
rect 13721 21450 13787 21453
rect 22510 21450 22570 21526
rect 27889 21523 27955 21526
rect 22829 21452 22895 21453
rect 22829 21450 22876 21452
rect 13721 21448 22570 21450
rect 13721 21392 13726 21448
rect 13782 21392 22570 21448
rect 13721 21390 22570 21392
rect 22784 21448 22876 21450
rect 22784 21392 22834 21448
rect 22784 21390 22876 21392
rect 13721 21387 13787 21390
rect 22829 21388 22876 21390
rect 22940 21388 22946 21452
rect 27705 21450 27771 21453
rect 36813 21450 36879 21453
rect 27705 21448 36879 21450
rect 27705 21392 27710 21448
rect 27766 21392 36818 21448
rect 36874 21392 36879 21448
rect 27705 21390 36879 21392
rect 22829 21387 22895 21388
rect 27705 21387 27771 21390
rect 36813 21387 36879 21390
rect 10041 21314 10107 21317
rect 20989 21314 21055 21317
rect 10041 21312 21055 21314
rect 10041 21256 10046 21312
rect 10102 21256 20994 21312
rect 21050 21256 21055 21312
rect 10041 21254 21055 21256
rect 10041 21251 10107 21254
rect 20989 21251 21055 21254
rect 22921 21314 22987 21317
rect 26049 21314 26115 21317
rect 22921 21312 26115 21314
rect 22921 21256 22926 21312
rect 22982 21256 26054 21312
rect 26110 21256 26115 21312
rect 22921 21254 26115 21256
rect 22921 21251 22987 21254
rect 26049 21251 26115 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 5717 21178 5783 21181
rect 24853 21178 24919 21181
rect 5717 21176 24919 21178
rect 5717 21120 5722 21176
rect 5778 21120 24858 21176
rect 24914 21120 24919 21176
rect 5717 21118 24919 21120
rect 5717 21115 5783 21118
rect 24853 21115 24919 21118
rect 25037 21178 25103 21181
rect 27705 21178 27771 21181
rect 25037 21176 27771 21178
rect 25037 21120 25042 21176
rect 25098 21120 27710 21176
rect 27766 21120 27771 21176
rect 25037 21118 27771 21120
rect 25037 21115 25103 21118
rect 27705 21115 27771 21118
rect 14181 21044 14247 21045
rect 14181 21042 14228 21044
rect 14136 21040 14228 21042
rect 14136 20984 14186 21040
rect 14136 20982 14228 20984
rect 14181 20980 14228 20982
rect 14292 20980 14298 21044
rect 14181 20979 14247 20980
rect 5625 20906 5691 20909
rect 22369 20906 22435 20909
rect 5625 20904 22435 20906
rect 5625 20848 5630 20904
rect 5686 20848 22374 20904
rect 22430 20848 22435 20904
rect 5625 20846 22435 20848
rect 5625 20843 5691 20846
rect 22369 20843 22435 20846
rect 9581 20772 9647 20773
rect 9581 20768 9628 20772
rect 9692 20770 9698 20772
rect 20345 20770 20411 20773
rect 21817 20770 21883 20773
rect 9581 20712 9586 20768
rect 9581 20708 9628 20712
rect 9692 20710 9738 20770
rect 20345 20768 21883 20770
rect 20345 20712 20350 20768
rect 20406 20712 21822 20768
rect 21878 20712 21883 20768
rect 20345 20710 21883 20712
rect 9692 20708 9698 20710
rect 9581 20707 9647 20708
rect 20345 20707 20411 20710
rect 21817 20707 21883 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 1485 20634 1551 20637
rect 798 20632 1551 20634
rect 798 20576 1490 20632
rect 1546 20576 1551 20632
rect 798 20574 1551 20576
rect 798 20528 858 20574
rect 1485 20571 1551 20574
rect 18137 20634 18203 20637
rect 19057 20634 19123 20637
rect 18137 20632 19123 20634
rect 18137 20576 18142 20632
rect 18198 20576 19062 20632
rect 19118 20576 19123 20632
rect 18137 20574 19123 20576
rect 18137 20571 18203 20574
rect 19057 20571 19123 20574
rect 25313 20634 25379 20637
rect 25446 20634 25452 20636
rect 25313 20632 25452 20634
rect 25313 20576 25318 20632
rect 25374 20576 25452 20632
rect 25313 20574 25452 20576
rect 25313 20571 25379 20574
rect 25446 20572 25452 20574
rect 25516 20572 25522 20636
rect 0 20438 858 20528
rect 10133 20498 10199 20501
rect 21909 20498 21975 20501
rect 10133 20496 21975 20498
rect 10133 20440 10138 20496
rect 10194 20440 21914 20496
rect 21970 20440 21975 20496
rect 10133 20438 21975 20440
rect 0 20408 800 20438
rect 10133 20435 10199 20438
rect 21909 20435 21975 20438
rect 38377 20498 38443 20501
rect 38618 20498 39418 20528
rect 38377 20496 39418 20498
rect 38377 20440 38382 20496
rect 38438 20440 39418 20496
rect 38377 20438 39418 20440
rect 38377 20435 38443 20438
rect 38618 20408 39418 20438
rect 9029 20362 9095 20365
rect 22369 20364 22435 20365
rect 22318 20362 22324 20364
rect 9029 20360 22324 20362
rect 22388 20362 22435 20364
rect 22388 20360 22516 20362
rect 9029 20304 9034 20360
rect 9090 20304 22324 20360
rect 22430 20304 22516 20360
rect 9029 20302 22324 20304
rect 9029 20299 9095 20302
rect 22318 20300 22324 20302
rect 22388 20302 22516 20304
rect 22388 20300 22435 20302
rect 22369 20299 22435 20300
rect 8569 20226 8635 20229
rect 23381 20226 23447 20229
rect 8569 20224 23447 20226
rect 8569 20168 8574 20224
rect 8630 20168 23386 20224
rect 23442 20168 23447 20224
rect 8569 20166 23447 20168
rect 8569 20163 8635 20166
rect 23381 20163 23447 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 17217 20090 17283 20093
rect 26049 20090 26115 20093
rect 17217 20088 26115 20090
rect 17217 20032 17222 20088
rect 17278 20032 26054 20088
rect 26110 20032 26115 20088
rect 17217 20030 26115 20032
rect 17217 20027 17283 20030
rect 26049 20027 26115 20030
rect 9489 19954 9555 19957
rect 22093 19954 22159 19957
rect 27337 19954 27403 19957
rect 9489 19952 27403 19954
rect 9489 19896 9494 19952
rect 9550 19896 22098 19952
rect 22154 19896 27342 19952
rect 27398 19896 27403 19952
rect 9489 19894 27403 19896
rect 9489 19891 9555 19894
rect 22093 19891 22159 19894
rect 27337 19891 27403 19894
rect 28993 19954 29059 19957
rect 30649 19954 30715 19957
rect 28993 19952 30715 19954
rect 28993 19896 28998 19952
rect 29054 19896 30654 19952
rect 30710 19896 30715 19952
rect 28993 19894 30715 19896
rect 28993 19891 29059 19894
rect 30649 19891 30715 19894
rect 8385 19818 8451 19821
rect 17217 19818 17283 19821
rect 23473 19818 23539 19821
rect 8385 19816 17283 19818
rect 8385 19760 8390 19816
rect 8446 19760 17222 19816
rect 17278 19760 17283 19816
rect 8385 19758 17283 19760
rect 8385 19755 8451 19758
rect 17217 19755 17283 19758
rect 19290 19816 23539 19818
rect 19290 19760 23478 19816
rect 23534 19760 23539 19816
rect 19290 19758 23539 19760
rect 12893 19682 12959 19685
rect 19290 19682 19350 19758
rect 23473 19755 23539 19758
rect 24025 19818 24091 19821
rect 26325 19818 26391 19821
rect 24025 19816 26391 19818
rect 24025 19760 24030 19816
rect 24086 19760 26330 19816
rect 26386 19760 26391 19816
rect 24025 19758 26391 19760
rect 24025 19755 24091 19758
rect 26325 19755 26391 19758
rect 12893 19680 19350 19682
rect 12893 19624 12898 19680
rect 12954 19624 19350 19680
rect 12893 19622 19350 19624
rect 23381 19682 23447 19685
rect 29085 19682 29151 19685
rect 23381 19680 29151 19682
rect 23381 19624 23386 19680
rect 23442 19624 29090 19680
rect 29146 19624 29151 19680
rect 23381 19622 29151 19624
rect 12893 19619 12959 19622
rect 23381 19619 23447 19622
rect 29085 19619 29151 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 13721 19546 13787 19549
rect 14641 19546 14707 19549
rect 13721 19544 14707 19546
rect 13721 19488 13726 19544
rect 13782 19488 14646 19544
rect 14702 19488 14707 19544
rect 13721 19486 14707 19488
rect 13721 19483 13787 19486
rect 14641 19483 14707 19486
rect 22369 19546 22435 19549
rect 25773 19546 25839 19549
rect 27613 19546 27679 19549
rect 22369 19544 27679 19546
rect 22369 19488 22374 19544
rect 22430 19488 25778 19544
rect 25834 19488 27618 19544
rect 27674 19488 27679 19544
rect 22369 19486 27679 19488
rect 22369 19483 22435 19486
rect 25773 19483 25839 19486
rect 27613 19483 27679 19486
rect 7925 19410 7991 19413
rect 25313 19410 25379 19413
rect 7925 19408 25379 19410
rect 7925 19352 7930 19408
rect 7986 19352 25318 19408
rect 25374 19352 25379 19408
rect 7925 19350 25379 19352
rect 7925 19347 7991 19350
rect 25313 19347 25379 19350
rect 27061 19410 27127 19413
rect 27889 19410 27955 19413
rect 27061 19408 27955 19410
rect 27061 19352 27066 19408
rect 27122 19352 27894 19408
rect 27950 19352 27955 19408
rect 27061 19350 27955 19352
rect 27061 19347 27127 19350
rect 27889 19347 27955 19350
rect 28257 19410 28323 19413
rect 31109 19410 31175 19413
rect 28257 19408 31175 19410
rect 28257 19352 28262 19408
rect 28318 19352 31114 19408
rect 31170 19352 31175 19408
rect 28257 19350 31175 19352
rect 28257 19347 28323 19350
rect 31109 19347 31175 19350
rect 22093 19274 22159 19277
rect 24301 19274 24367 19277
rect 22093 19272 24367 19274
rect 22093 19216 22098 19272
rect 22154 19216 24306 19272
rect 24362 19216 24367 19272
rect 22093 19214 24367 19216
rect 22093 19211 22159 19214
rect 24301 19211 24367 19214
rect 11237 19138 11303 19141
rect 24945 19138 25011 19141
rect 11237 19136 25011 19138
rect 11237 19080 11242 19136
rect 11298 19080 24950 19136
rect 25006 19080 25011 19136
rect 11237 19078 25011 19080
rect 11237 19075 11303 19078
rect 24945 19075 25011 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 15694 18940 15700 19004
rect 15764 19002 15770 19004
rect 22369 19002 22435 19005
rect 15764 19000 22435 19002
rect 15764 18944 22374 19000
rect 22430 18944 22435 19000
rect 15764 18942 22435 18944
rect 15764 18940 15770 18942
rect 22369 18939 22435 18942
rect 5993 18866 6059 18869
rect 23565 18866 23631 18869
rect 5993 18864 23631 18866
rect 5993 18808 5998 18864
rect 6054 18808 23570 18864
rect 23626 18808 23631 18864
rect 5993 18806 23631 18808
rect 5993 18803 6059 18806
rect 23565 18803 23631 18806
rect 15653 18730 15719 18733
rect 18045 18730 18111 18733
rect 18413 18730 18479 18733
rect 15653 18728 18479 18730
rect 15653 18672 15658 18728
rect 15714 18672 18050 18728
rect 18106 18672 18418 18728
rect 18474 18672 18479 18728
rect 15653 18670 18479 18672
rect 15653 18667 15719 18670
rect 18045 18667 18111 18670
rect 18413 18667 18479 18670
rect 19570 18528 19886 18529
rect 0 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 14733 18322 14799 18325
rect 19057 18322 19123 18325
rect 14733 18320 19123 18322
rect 14733 18264 14738 18320
rect 14794 18264 19062 18320
rect 19118 18264 19123 18320
rect 14733 18262 19123 18264
rect 14733 18259 14799 18262
rect 19057 18259 19123 18262
rect 30373 18322 30439 18325
rect 33777 18322 33843 18325
rect 30373 18320 33843 18322
rect 30373 18264 30378 18320
rect 30434 18264 33782 18320
rect 33838 18264 33843 18320
rect 30373 18262 33843 18264
rect 30373 18259 30439 18262
rect 33777 18259 33843 18262
rect 18229 18186 18295 18189
rect 18965 18186 19031 18189
rect 18229 18184 19031 18186
rect 18229 18128 18234 18184
rect 18290 18128 18970 18184
rect 19026 18128 19031 18184
rect 18229 18126 19031 18128
rect 18229 18123 18295 18126
rect 18965 18123 19031 18126
rect 10869 18050 10935 18053
rect 10869 18048 17234 18050
rect 10869 17992 10874 18048
rect 10930 17992 17234 18048
rect 10869 17990 17234 17992
rect 10869 17987 10935 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 9029 17914 9095 17917
rect 9806 17914 9812 17916
rect 9029 17912 9812 17914
rect 9029 17856 9034 17912
rect 9090 17856 9812 17912
rect 9029 17854 9812 17856
rect 9029 17851 9095 17854
rect 9806 17852 9812 17854
rect 9876 17852 9882 17916
rect 17174 17778 17234 17990
rect 20110 17988 20116 18052
rect 20180 18050 20186 18052
rect 21449 18050 21515 18053
rect 20180 18048 21515 18050
rect 20180 17992 21454 18048
rect 21510 17992 21515 18048
rect 20180 17990 21515 17992
rect 20180 17988 20186 17990
rect 21449 17987 21515 17990
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 17534 17852 17540 17916
rect 17604 17914 17610 17916
rect 18229 17914 18295 17917
rect 17604 17912 18295 17914
rect 17604 17856 18234 17912
rect 18290 17856 18295 17912
rect 17604 17854 18295 17856
rect 17604 17852 17610 17854
rect 18229 17851 18295 17854
rect 18413 17916 18479 17917
rect 18413 17912 18460 17916
rect 18524 17914 18530 17916
rect 18413 17856 18418 17912
rect 18413 17852 18460 17856
rect 18524 17854 18570 17914
rect 18524 17852 18530 17854
rect 21950 17852 21956 17916
rect 22020 17914 22026 17916
rect 22645 17914 22711 17917
rect 22020 17912 22711 17914
rect 22020 17856 22650 17912
rect 22706 17856 22711 17912
rect 22020 17854 22711 17856
rect 22020 17852 22026 17854
rect 18413 17851 18479 17852
rect 22645 17851 22711 17854
rect 23381 17914 23447 17917
rect 23606 17914 23612 17916
rect 23381 17912 23612 17914
rect 23381 17856 23386 17912
rect 23442 17856 23612 17912
rect 23381 17854 23612 17856
rect 23381 17851 23447 17854
rect 23606 17852 23612 17854
rect 23676 17852 23682 17916
rect 27705 17778 27771 17781
rect 17174 17776 27771 17778
rect 17174 17720 27710 17776
rect 27766 17720 27771 17776
rect 17174 17718 27771 17720
rect 27705 17715 27771 17718
rect 38377 17778 38443 17781
rect 38618 17778 39418 17808
rect 38377 17776 39418 17778
rect 38377 17720 38382 17776
rect 38438 17720 39418 17776
rect 38377 17718 39418 17720
rect 38377 17715 38443 17718
rect 38618 17688 39418 17718
rect 23197 17642 23263 17645
rect 26182 17642 26188 17644
rect 23197 17640 26188 17642
rect 23197 17584 23202 17640
rect 23258 17584 26188 17640
rect 23197 17582 26188 17584
rect 23197 17579 23263 17582
rect 26182 17580 26188 17582
rect 26252 17580 26258 17644
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 32029 17234 32095 17237
rect 32857 17234 32923 17237
rect 32029 17232 32923 17234
rect 32029 17176 32034 17232
rect 32090 17176 32862 17232
rect 32918 17176 32923 17232
rect 32029 17174 32923 17176
rect 32029 17171 32095 17174
rect 32857 17171 32923 17174
rect 24669 17100 24735 17101
rect 24669 17098 24716 17100
rect 24624 17096 24716 17098
rect 24624 17040 24674 17096
rect 24624 17038 24716 17040
rect 24669 17036 24716 17038
rect 24780 17036 24786 17100
rect 24669 17035 24735 17036
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19333 16554 19399 16557
rect 23289 16554 23355 16557
rect 24485 16556 24551 16557
rect 24485 16554 24532 16556
rect 19333 16552 23355 16554
rect 19333 16496 19338 16552
rect 19394 16496 23294 16552
rect 23350 16496 23355 16552
rect 19333 16494 23355 16496
rect 24440 16552 24532 16554
rect 24440 16496 24490 16552
rect 24440 16494 24532 16496
rect 19333 16491 19399 16494
rect 23289 16491 23355 16494
rect 24485 16492 24532 16494
rect 24596 16492 24602 16556
rect 24485 16491 24551 16492
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 12341 16146 12407 16149
rect 24485 16146 24551 16149
rect 12341 16144 24551 16146
rect 12341 16088 12346 16144
rect 12402 16088 24490 16144
rect 24546 16088 24551 16144
rect 12341 16086 24551 16088
rect 12341 16083 12407 16086
rect 24485 16083 24551 16086
rect 29177 16146 29243 16149
rect 29637 16146 29703 16149
rect 29177 16144 29703 16146
rect 29177 16088 29182 16144
rect 29238 16088 29642 16144
rect 29698 16088 29703 16144
rect 29177 16086 29703 16088
rect 29177 16083 29243 16086
rect 29637 16083 29703 16086
rect 12249 16010 12315 16013
rect 23749 16010 23815 16013
rect 12249 16008 23815 16010
rect 12249 15952 12254 16008
rect 12310 15952 23754 16008
rect 23810 15952 23815 16008
rect 12249 15950 23815 15952
rect 12249 15947 12315 15950
rect 23749 15947 23815 15950
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 933 15738 999 15741
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 37825 15738 37891 15741
rect 38618 15738 39418 15768
rect 37825 15736 39418 15738
rect 37825 15680 37830 15736
rect 37886 15680 39418 15736
rect 37825 15678 39418 15680
rect 37825 15675 37891 15678
rect 38618 15648 39418 15678
rect 11329 15602 11395 15605
rect 17585 15602 17651 15605
rect 11329 15600 17651 15602
rect 11329 15544 11334 15600
rect 11390 15544 17590 15600
rect 17646 15544 17651 15600
rect 11329 15542 17651 15544
rect 11329 15539 11395 15542
rect 17585 15539 17651 15542
rect 11513 15466 11579 15469
rect 25129 15466 25195 15469
rect 11513 15464 25195 15466
rect 11513 15408 11518 15464
rect 11574 15408 25134 15464
rect 25190 15408 25195 15464
rect 11513 15406 25195 15408
rect 11513 15403 11579 15406
rect 25129 15403 25195 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 27613 15194 27679 15197
rect 28441 15194 28507 15197
rect 27613 15192 28507 15194
rect 27613 15136 27618 15192
rect 27674 15136 28446 15192
rect 28502 15136 28507 15192
rect 27613 15134 28507 15136
rect 27613 15131 27679 15134
rect 28441 15131 28507 15134
rect 23197 15058 23263 15061
rect 28717 15058 28783 15061
rect 23197 15056 28783 15058
rect 23197 15000 23202 15056
rect 23258 15000 28722 15056
rect 28778 15000 28783 15056
rect 23197 14998 28783 15000
rect 23197 14995 23263 14998
rect 28717 14995 28783 14998
rect 26325 14922 26391 14925
rect 28533 14922 28599 14925
rect 26325 14920 28599 14922
rect 26325 14864 26330 14920
rect 26386 14864 28538 14920
rect 28594 14864 28599 14920
rect 26325 14862 28599 14864
rect 26325 14859 26391 14862
rect 28533 14859 28599 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 14365 14514 14431 14517
rect 17769 14514 17835 14517
rect 14365 14512 17835 14514
rect 14365 14456 14370 14512
rect 14426 14456 17774 14512
rect 17830 14456 17835 14512
rect 14365 14454 17835 14456
rect 14365 14451 14431 14454
rect 17769 14451 17835 14454
rect 9581 14378 9647 14381
rect 30189 14378 30255 14381
rect 9581 14376 30255 14378
rect 9581 14320 9586 14376
rect 9642 14320 30194 14376
rect 30250 14320 30255 14376
rect 9581 14318 30255 14320
rect 9581 14315 9647 14318
rect 30189 14315 30255 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 9581 13700 9647 13701
rect 9581 13698 9628 13700
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 9536 13696 9628 13698
rect 9536 13640 9586 13696
rect 9536 13638 9628 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 9581 13636 9628 13638
rect 9692 13636 9698 13700
rect 9581 13635 9647 13636
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 38618 13608 39418 13728
rect 34930 13567 35246 13568
rect 26734 13364 26740 13428
rect 26804 13426 26810 13428
rect 27613 13426 27679 13429
rect 26804 13424 27679 13426
rect 26804 13368 27618 13424
rect 27674 13368 27679 13424
rect 26804 13366 27679 13368
rect 26804 13364 26810 13366
rect 27613 13363 27679 13366
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 10225 13018 10291 13021
rect 18689 13018 18755 13021
rect 10225 13016 18755 13018
rect 10225 12960 10230 13016
rect 10286 12960 18694 13016
rect 18750 12960 18755 13016
rect 10225 12958 18755 12960
rect 10225 12955 10291 12958
rect 18689 12955 18755 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 18689 11658 18755 11661
rect 27705 11658 27771 11661
rect 18689 11656 27771 11658
rect 18689 11600 18694 11656
rect 18750 11600 27710 11656
rect 27766 11600 27771 11656
rect 18689 11598 27771 11600
rect 18689 11595 18755 11598
rect 27705 11595 27771 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 21449 10978 21515 10981
rect 22553 10978 22619 10981
rect 21449 10976 22619 10978
rect 21449 10920 21454 10976
rect 21510 10920 22558 10976
rect 22614 10920 22619 10976
rect 21449 10918 22619 10920
rect 21449 10915 21515 10918
rect 22553 10915 22619 10918
rect 37917 10978 37983 10981
rect 38618 10978 39418 11008
rect 37917 10976 39418 10978
rect 37917 10920 37922 10976
rect 37978 10920 39418 10976
rect 37917 10918 39418 10920
rect 37917 10915 37983 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 38618 10888 39418 10918
rect 19570 10847 19886 10848
rect 21541 10706 21607 10709
rect 23013 10706 23079 10709
rect 21541 10704 23079 10706
rect 21541 10648 21546 10704
rect 21602 10648 23018 10704
rect 23074 10648 23079 10704
rect 21541 10646 23079 10648
rect 21541 10643 21607 10646
rect 23013 10643 23079 10646
rect 17493 10570 17559 10573
rect 27889 10570 27955 10573
rect 17493 10568 27955 10570
rect 17493 10512 17498 10568
rect 17554 10512 27894 10568
rect 27950 10512 27955 10568
rect 17493 10510 27955 10512
rect 17493 10507 17559 10510
rect 27889 10507 27955 10510
rect 16430 10372 16436 10436
rect 16500 10434 16506 10436
rect 18229 10434 18295 10437
rect 16500 10432 18295 10434
rect 16500 10376 18234 10432
rect 18290 10376 18295 10432
rect 16500 10374 18295 10376
rect 16500 10372 16506 10374
rect 18229 10371 18295 10374
rect 20805 10434 20871 10437
rect 27981 10434 28047 10437
rect 28625 10434 28691 10437
rect 20805 10432 28691 10434
rect 20805 10376 20810 10432
rect 20866 10376 27986 10432
rect 28042 10376 28630 10432
rect 28686 10376 28691 10432
rect 20805 10374 28691 10376
rect 20805 10371 20871 10374
rect 27981 10371 28047 10374
rect 28625 10371 28691 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 30189 10162 30255 10165
rect 32857 10162 32923 10165
rect 30189 10160 32923 10162
rect 30189 10104 30194 10160
rect 30250 10104 32862 10160
rect 32918 10104 32923 10160
rect 30189 10102 32923 10104
rect 30189 10099 30255 10102
rect 32857 10099 32923 10102
rect 20345 9890 20411 9893
rect 24117 9890 24183 9893
rect 24485 9890 24551 9893
rect 20345 9888 24551 9890
rect 20345 9832 20350 9888
rect 20406 9832 24122 9888
rect 24178 9832 24490 9888
rect 24546 9832 24551 9888
rect 20345 9830 24551 9832
rect 20345 9827 20411 9830
rect 24117 9827 24183 9830
rect 24485 9827 24551 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 3233 9618 3299 9621
rect 22277 9620 22343 9621
rect 22277 9618 22324 9620
rect 3233 9616 22110 9618
rect 3233 9560 3238 9616
rect 3294 9560 22110 9616
rect 3233 9558 22110 9560
rect 22232 9616 22324 9618
rect 22232 9560 22282 9616
rect 22232 9558 22324 9560
rect 3233 9555 3299 9558
rect 22050 9482 22110 9558
rect 22277 9556 22324 9558
rect 22388 9556 22394 9620
rect 22277 9555 22343 9556
rect 30005 9482 30071 9485
rect 30649 9482 30715 9485
rect 22050 9480 30715 9482
rect 22050 9424 30010 9480
rect 30066 9424 30654 9480
rect 30710 9424 30715 9480
rect 22050 9422 30715 9424
rect 30005 9419 30071 9422
rect 30649 9419 30715 9422
rect 23749 9346 23815 9349
rect 24761 9346 24827 9349
rect 23749 9344 24827 9346
rect 23749 9288 23754 9344
rect 23810 9288 24766 9344
rect 24822 9288 24827 9344
rect 23749 9286 24827 9288
rect 23749 9283 23815 9286
rect 24761 9283 24827 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 23933 9210 23999 9213
rect 25497 9210 25563 9213
rect 23933 9208 25563 9210
rect 23933 9152 23938 9208
rect 23994 9152 25502 9208
rect 25558 9152 25563 9208
rect 23933 9150 25563 9152
rect 23933 9147 23999 9150
rect 25497 9147 25563 9150
rect 4153 9074 4219 9077
rect 22829 9074 22895 9077
rect 24710 9074 24716 9076
rect 4153 9072 24716 9074
rect 4153 9016 4158 9072
rect 4214 9016 22834 9072
rect 22890 9016 24716 9072
rect 4153 9014 24716 9016
rect 4153 9011 4219 9014
rect 22829 9011 22895 9014
rect 24710 9012 24716 9014
rect 24780 9012 24786 9076
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 26877 8938 26943 8941
rect 27981 8938 28047 8941
rect 26877 8936 28047 8938
rect 26877 8880 26882 8936
rect 26938 8880 27986 8936
rect 28042 8880 28047 8936
rect 26877 8878 28047 8880
rect 26877 8875 26943 8878
rect 27981 8875 28047 8878
rect 38285 8938 38351 8941
rect 38618 8938 39418 8968
rect 38285 8936 39418 8938
rect 38285 8880 38290 8936
rect 38346 8880 39418 8936
rect 38285 8878 39418 8880
rect 38285 8875 38351 8878
rect 38618 8848 39418 8878
rect 26325 8802 26391 8805
rect 27797 8802 27863 8805
rect 26325 8800 27863 8802
rect 26325 8744 26330 8800
rect 26386 8744 27802 8800
rect 27858 8744 27863 8800
rect 26325 8742 27863 8744
rect 26325 8739 26391 8742
rect 27797 8739 27863 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 12157 8530 12223 8533
rect 14917 8530 14983 8533
rect 18965 8532 19031 8533
rect 18965 8530 19012 8532
rect 12157 8528 14983 8530
rect 12157 8472 12162 8528
rect 12218 8472 14922 8528
rect 14978 8472 14983 8528
rect 12157 8470 14983 8472
rect 18920 8528 19012 8530
rect 18920 8472 18970 8528
rect 18920 8470 19012 8472
rect 12157 8467 12223 8470
rect 14917 8467 14983 8470
rect 18965 8468 19012 8470
rect 19076 8468 19082 8532
rect 18965 8467 19031 8468
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 18229 6900 18295 6901
rect 18229 6898 18276 6900
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 18184 6896 18276 6898
rect 18184 6840 18234 6896
rect 18184 6838 18276 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 18229 6836 18276 6838
rect 18340 6836 18346 6900
rect 18229 6835 18295 6836
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 38618 6128 39418 6248
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 21817 4586 21883 4589
rect 25129 4586 25195 4589
rect 25589 4586 25655 4589
rect 21817 4584 25655 4586
rect 21817 4528 21822 4584
rect 21878 4528 25134 4584
rect 25190 4528 25594 4584
rect 25650 4528 25655 4584
rect 21817 4526 25655 4528
rect 21817 4523 21883 4526
rect 25129 4523 25195 4526
rect 25589 4523 25655 4526
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 38618 4088 39418 4208
rect 12525 4044 12591 4045
rect 12525 4040 12572 4044
rect 12636 4042 12642 4044
rect 13169 4042 13235 4045
rect 13302 4042 13308 4044
rect 12525 3984 12530 4040
rect 12525 3980 12572 3984
rect 12636 3982 12682 4042
rect 13169 4040 13308 4042
rect 13169 3984 13174 4040
rect 13230 3984 13308 4040
rect 13169 3982 13308 3984
rect 12636 3980 12642 3982
rect 12525 3979 12591 3980
rect 13169 3979 13235 3982
rect 13302 3980 13308 3982
rect 13372 3980 13378 4044
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 0 2048 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 37181 1458 37247 1461
rect 38618 1458 39418 1488
rect 37181 1456 39418 1458
rect 37181 1400 37186 1456
rect 37242 1400 39418 1456
rect 37181 1398 39418 1400
rect 37181 1395 37247 1398
rect 38618 1368 39418 1398
<< via3 >>
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 14228 38932 14292 38996
rect 9812 38796 9876 38860
rect 10364 38660 10428 38724
rect 22876 38660 22940 38724
rect 23980 38660 24044 38724
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 22140 37300 22204 37364
rect 25268 37360 25332 37364
rect 25268 37304 25282 37360
rect 25282 37304 25332 37360
rect 25268 37300 25332 37304
rect 27844 37300 27908 37364
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 17540 35940 17604 36004
rect 20300 35940 20364 36004
rect 20484 36000 20548 36004
rect 20484 35944 20498 36000
rect 20498 35944 20548 36000
rect 20484 35940 20548 35944
rect 28948 35940 29012 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 14780 35668 14844 35732
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 26188 33900 26252 33964
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 21220 33492 21284 33556
rect 19012 33280 19076 33284
rect 19012 33224 19062 33280
rect 19062 33224 19076 33280
rect 19012 33220 19076 33224
rect 24532 33220 24596 33284
rect 25452 33280 25516 33284
rect 25452 33224 25466 33280
rect 25466 33224 25516 33280
rect 25452 33220 25516 33224
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 28948 33084 29012 33148
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 18092 32132 18156 32196
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 15700 31996 15764 32060
rect 18276 31996 18340 32060
rect 28948 31996 29012 32060
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 21220 31316 21284 31380
rect 27844 31044 27908 31108
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 18460 30364 18524 30428
rect 23980 30364 24044 30428
rect 26740 30424 26804 30428
rect 26740 30368 26754 30424
rect 26754 30368 26804 30424
rect 26740 30364 26804 30368
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 21220 29412 21284 29476
rect 13308 29004 13372 29068
rect 16436 29004 16500 29068
rect 23612 29064 23676 29068
rect 23612 29008 23626 29064
rect 23626 29008 23676 29064
rect 23612 29004 23676 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 18092 28792 18156 28796
rect 18092 28736 18106 28792
rect 18106 28736 18156 28792
rect 18092 28732 18156 28736
rect 20300 28656 20364 28660
rect 20300 28600 20314 28656
rect 20314 28600 20364 28656
rect 20300 28596 20364 28600
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 25820 28188 25884 28252
rect 28948 27916 29012 27980
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 21956 27704 22020 27708
rect 21956 27648 21970 27704
rect 21970 27648 22020 27704
rect 21956 27644 22020 27648
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 20116 26344 20180 26348
rect 20116 26288 20130 26344
rect 20130 26288 20180 26344
rect 20116 26284 20180 26288
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 25268 26012 25332 26076
rect 20484 25740 20548 25804
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 22140 24168 22204 24172
rect 22140 24112 22154 24168
rect 22154 24112 22204 24168
rect 22140 24108 22204 24112
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 25820 23760 25884 23764
rect 25820 23704 25870 23760
rect 25870 23704 25884 23760
rect 25820 23700 25884 23704
rect 12572 23488 12636 23492
rect 12572 23432 12622 23488
rect 12622 23432 12636 23488
rect 12572 23428 12636 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 14780 21720 14844 21724
rect 14780 21664 14794 21720
rect 14794 21664 14844 21720
rect 14780 21660 14844 21664
rect 9812 21524 9876 21588
rect 10364 21584 10428 21588
rect 10364 21528 10378 21584
rect 10378 21528 10428 21584
rect 10364 21524 10428 21528
rect 22876 21448 22940 21452
rect 22876 21392 22890 21448
rect 22890 21392 22940 21448
rect 22876 21388 22940 21392
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 14228 21040 14292 21044
rect 14228 20984 14242 21040
rect 14242 20984 14292 21040
rect 14228 20980 14292 20984
rect 9628 20768 9692 20772
rect 9628 20712 9642 20768
rect 9642 20712 9692 20768
rect 9628 20708 9692 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 25452 20572 25516 20636
rect 22324 20360 22388 20364
rect 22324 20304 22374 20360
rect 22374 20304 22388 20360
rect 22324 20300 22388 20304
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 15700 18940 15764 19004
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 9812 17852 9876 17916
rect 20116 17988 20180 18052
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 17540 17852 17604 17916
rect 18460 17912 18524 17916
rect 18460 17856 18474 17912
rect 18474 17856 18524 17912
rect 18460 17852 18524 17856
rect 21956 17852 22020 17916
rect 23612 17852 23676 17916
rect 26188 17580 26252 17644
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 24716 17096 24780 17100
rect 24716 17040 24730 17096
rect 24730 17040 24780 17096
rect 24716 17036 24780 17040
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 24532 16552 24596 16556
rect 24532 16496 24546 16552
rect 24546 16496 24596 16552
rect 24532 16492 24596 16496
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 9628 13696 9692 13700
rect 9628 13640 9642 13696
rect 9642 13640 9692 13696
rect 9628 13636 9692 13640
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 26740 13364 26804 13428
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 16436 10372 16500 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 22324 9616 22388 9620
rect 22324 9560 22338 9616
rect 22338 9560 22388 9616
rect 22324 9556 22388 9560
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 24716 9012 24780 9076
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 19012 8528 19076 8532
rect 19012 8472 19026 8528
rect 19026 8472 19076 8528
rect 19012 8468 19076 8472
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 18276 6896 18340 6900
rect 18276 6840 18290 6896
rect 18290 6840 18340 6896
rect 18276 6836 18340 6840
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 12572 4040 12636 4044
rect 12572 3984 12586 4040
rect 12586 3984 12636 4040
rect 12572 3980 12636 3984
rect 13308 3980 13372 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 38656 4528 39216
rect 19568 39200 19888 39216
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 14227 38996 14293 38997
rect 14227 38932 14228 38996
rect 14292 38932 14293 38996
rect 14227 38931 14293 38932
rect 9811 38860 9877 38861
rect 9811 38796 9812 38860
rect 9876 38796 9877 38860
rect 9811 38795 9877 38796
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 9814 21589 9874 38795
rect 10363 38724 10429 38725
rect 10363 38660 10364 38724
rect 10428 38660 10429 38724
rect 10363 38659 10429 38660
rect 10366 21589 10426 38659
rect 13307 29068 13373 29069
rect 13307 29004 13308 29068
rect 13372 29004 13373 29068
rect 13307 29003 13373 29004
rect 12571 23492 12637 23493
rect 12571 23428 12572 23492
rect 12636 23428 12637 23492
rect 12571 23427 12637 23428
rect 9811 21588 9877 21589
rect 9811 21524 9812 21588
rect 9876 21524 9877 21588
rect 9811 21523 9877 21524
rect 10363 21588 10429 21589
rect 10363 21524 10364 21588
rect 10428 21524 10429 21588
rect 10363 21523 10429 21524
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 9627 20772 9693 20773
rect 9627 20708 9628 20772
rect 9692 20708 9693 20772
rect 9627 20707 9693 20708
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 9630 13701 9690 20707
rect 9814 17917 9874 21523
rect 9811 17916 9877 17917
rect 9811 17852 9812 17916
rect 9876 17852 9877 17916
rect 9811 17851 9877 17852
rect 9627 13700 9693 13701
rect 9627 13636 9628 13700
rect 9692 13636 9693 13700
rect 9627 13635 9693 13636
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 12574 4045 12634 23427
rect 13310 4045 13370 29003
rect 14230 21045 14290 38931
rect 19568 38112 19888 39136
rect 22875 38724 22941 38725
rect 22875 38660 22876 38724
rect 22940 38660 22941 38724
rect 22875 38659 22941 38660
rect 23979 38724 24045 38725
rect 23979 38660 23980 38724
rect 24044 38660 24045 38724
rect 23979 38659 24045 38660
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 22139 37364 22205 37365
rect 22139 37300 22140 37364
rect 22204 37300 22205 37364
rect 22139 37299 22205 37300
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 17539 36004 17605 36005
rect 17539 35940 17540 36004
rect 17604 35940 17605 36004
rect 17539 35939 17605 35940
rect 14779 35732 14845 35733
rect 14779 35668 14780 35732
rect 14844 35668 14845 35732
rect 14779 35667 14845 35668
rect 14782 21725 14842 35667
rect 15699 32060 15765 32061
rect 15699 31996 15700 32060
rect 15764 31996 15765 32060
rect 15699 31995 15765 31996
rect 14779 21724 14845 21725
rect 14779 21660 14780 21724
rect 14844 21660 14845 21724
rect 14779 21659 14845 21660
rect 14227 21044 14293 21045
rect 14227 20980 14228 21044
rect 14292 20980 14293 21044
rect 14227 20979 14293 20980
rect 15702 19005 15762 31995
rect 16435 29068 16501 29069
rect 16435 29004 16436 29068
rect 16500 29004 16501 29068
rect 16435 29003 16501 29004
rect 15699 19004 15765 19005
rect 15699 18940 15700 19004
rect 15764 18940 15765 19004
rect 15699 18939 15765 18940
rect 16438 10437 16498 29003
rect 17542 17917 17602 35939
rect 19568 35936 19888 36960
rect 20299 36004 20365 36005
rect 20299 35940 20300 36004
rect 20364 35940 20365 36004
rect 20299 35939 20365 35940
rect 20483 36004 20549 36005
rect 20483 35940 20484 36004
rect 20548 35940 20549 36004
rect 20483 35939 20549 35940
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19011 33284 19077 33285
rect 19011 33220 19012 33284
rect 19076 33220 19077 33284
rect 19011 33219 19077 33220
rect 18091 32196 18157 32197
rect 18091 32132 18092 32196
rect 18156 32132 18157 32196
rect 18091 32131 18157 32132
rect 18094 28797 18154 32131
rect 18275 32060 18341 32061
rect 18275 31996 18276 32060
rect 18340 31996 18341 32060
rect 18275 31995 18341 31996
rect 18091 28796 18157 28797
rect 18091 28732 18092 28796
rect 18156 28732 18157 28796
rect 18091 28731 18157 28732
rect 17539 17916 17605 17917
rect 17539 17852 17540 17916
rect 17604 17852 17605 17916
rect 17539 17851 17605 17852
rect 16435 10436 16501 10437
rect 16435 10372 16436 10436
rect 16500 10372 16501 10436
rect 16435 10371 16501 10372
rect 18278 6901 18338 31995
rect 18459 30428 18525 30429
rect 18459 30364 18460 30428
rect 18524 30364 18525 30428
rect 18459 30363 18525 30364
rect 18462 17917 18522 30363
rect 18459 17916 18525 17917
rect 18459 17852 18460 17916
rect 18524 17852 18525 17916
rect 18459 17851 18525 17852
rect 19014 8533 19074 33219
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 20302 28661 20362 35939
rect 20299 28660 20365 28661
rect 20299 28596 20300 28660
rect 20364 28596 20365 28660
rect 20299 28595 20365 28596
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 20115 26348 20181 26349
rect 20115 26284 20116 26348
rect 20180 26284 20181 26348
rect 20115 26283 20181 26284
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 20118 18053 20178 26283
rect 20486 25805 20546 35939
rect 21219 33556 21285 33557
rect 21219 33492 21220 33556
rect 21284 33492 21285 33556
rect 21219 33491 21285 33492
rect 21222 31381 21282 33491
rect 21219 31380 21285 31381
rect 21219 31316 21220 31380
rect 21284 31316 21285 31380
rect 21219 31315 21285 31316
rect 21222 29477 21282 31315
rect 21219 29476 21285 29477
rect 21219 29412 21220 29476
rect 21284 29412 21285 29476
rect 21219 29411 21285 29412
rect 21955 27708 22021 27709
rect 21955 27644 21956 27708
rect 22020 27644 22021 27708
rect 21955 27643 22021 27644
rect 20483 25804 20549 25805
rect 20483 25740 20484 25804
rect 20548 25740 20549 25804
rect 20483 25739 20549 25740
rect 20115 18052 20181 18053
rect 20115 17988 20116 18052
rect 20180 17988 20181 18052
rect 20115 17987 20181 17988
rect 21958 17917 22018 27643
rect 22142 24173 22202 37299
rect 22139 24172 22205 24173
rect 22139 24108 22140 24172
rect 22204 24108 22205 24172
rect 22139 24107 22205 24108
rect 22878 21453 22938 38659
rect 23982 30429 24042 38659
rect 34928 38656 35248 39216
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 25267 37364 25333 37365
rect 25267 37300 25268 37364
rect 25332 37300 25333 37364
rect 25267 37299 25333 37300
rect 27843 37364 27909 37365
rect 27843 37300 27844 37364
rect 27908 37300 27909 37364
rect 27843 37299 27909 37300
rect 24531 33284 24597 33285
rect 24531 33220 24532 33284
rect 24596 33220 24597 33284
rect 24531 33219 24597 33220
rect 23979 30428 24045 30429
rect 23979 30364 23980 30428
rect 24044 30364 24045 30428
rect 23979 30363 24045 30364
rect 23611 29068 23677 29069
rect 23611 29004 23612 29068
rect 23676 29004 23677 29068
rect 23611 29003 23677 29004
rect 22875 21452 22941 21453
rect 22875 21388 22876 21452
rect 22940 21388 22941 21452
rect 22875 21387 22941 21388
rect 22323 20364 22389 20365
rect 22323 20300 22324 20364
rect 22388 20300 22389 20364
rect 22323 20299 22389 20300
rect 21955 17916 22021 17917
rect 21955 17852 21956 17916
rect 22020 17852 22021 17916
rect 21955 17851 22021 17852
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 22326 9621 22386 20299
rect 23614 17917 23674 29003
rect 23611 17916 23677 17917
rect 23611 17852 23612 17916
rect 23676 17852 23677 17916
rect 23611 17851 23677 17852
rect 24534 16557 24594 33219
rect 25270 26077 25330 37299
rect 26187 33964 26253 33965
rect 26187 33900 26188 33964
rect 26252 33900 26253 33964
rect 26187 33899 26253 33900
rect 25451 33284 25517 33285
rect 25451 33220 25452 33284
rect 25516 33220 25517 33284
rect 25451 33219 25517 33220
rect 25267 26076 25333 26077
rect 25267 26012 25268 26076
rect 25332 26012 25333 26076
rect 25267 26011 25333 26012
rect 25454 20637 25514 33219
rect 25819 28252 25885 28253
rect 25819 28188 25820 28252
rect 25884 28188 25885 28252
rect 25819 28187 25885 28188
rect 25822 23765 25882 28187
rect 25819 23764 25885 23765
rect 25819 23700 25820 23764
rect 25884 23700 25885 23764
rect 25819 23699 25885 23700
rect 25451 20636 25517 20637
rect 25451 20572 25452 20636
rect 25516 20572 25517 20636
rect 25451 20571 25517 20572
rect 26190 17645 26250 33899
rect 27846 31109 27906 37299
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 28947 36004 29013 36005
rect 28947 35940 28948 36004
rect 29012 35940 29013 36004
rect 28947 35939 29013 35940
rect 28950 33149 29010 35939
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 28947 33148 29013 33149
rect 28947 33084 28948 33148
rect 29012 33084 29013 33148
rect 28947 33083 29013 33084
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 28947 32060 29013 32061
rect 28947 31996 28948 32060
rect 29012 31996 29013 32060
rect 28947 31995 29013 31996
rect 27843 31108 27909 31109
rect 27843 31044 27844 31108
rect 27908 31044 27909 31108
rect 27843 31043 27909 31044
rect 26739 30428 26805 30429
rect 26739 30364 26740 30428
rect 26804 30364 26805 30428
rect 26739 30363 26805 30364
rect 26187 17644 26253 17645
rect 26187 17580 26188 17644
rect 26252 17580 26253 17644
rect 26187 17579 26253 17580
rect 24715 17100 24781 17101
rect 24715 17036 24716 17100
rect 24780 17036 24781 17100
rect 24715 17035 24781 17036
rect 24531 16556 24597 16557
rect 24531 16492 24532 16556
rect 24596 16492 24597 16556
rect 24531 16491 24597 16492
rect 22323 9620 22389 9621
rect 22323 9556 22324 9620
rect 22388 9556 22389 9620
rect 22323 9555 22389 9556
rect 24718 9077 24778 17035
rect 26742 13429 26802 30363
rect 28950 27981 29010 31995
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 28947 27980 29013 27981
rect 28947 27916 28948 27980
rect 29012 27916 29013 27980
rect 28947 27915 29013 27916
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 26739 13428 26805 13429
rect 26739 13364 26740 13428
rect 26804 13364 26805 13428
rect 26739 13363 26805 13364
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 24715 9076 24781 9077
rect 24715 9012 24716 9076
rect 24780 9012 24781 9076
rect 24715 9011 24781 9012
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19011 8532 19077 8533
rect 19011 8468 19012 8532
rect 19076 8468 19077 8532
rect 19011 8467 19077 8468
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 18275 6900 18341 6901
rect 18275 6836 18276 6900
rect 18340 6836 18341 6900
rect 18275 6835 18341 6836
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 12571 4044 12637 4045
rect 12571 3980 12572 4044
rect 12636 3980 12637 4044
rect 12571 3979 12637 3980
rect 13307 4044 13373 4045
rect 13307 3980 13308 4044
rect 13372 3980 13373 4044
rect 13307 3979 13373 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__inv_2  _1275_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20332 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _1276_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13156 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _1277_
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1278_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _1279_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1280_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13248 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1281_
timestamp 1688980957
transform 1 0 16836 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_1  _1282_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14996 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1283_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1284_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12696 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1285_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13984 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  _1286_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  _1287_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_2  _1288_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22172 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _1289_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15364 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__a21boi_1  _1290_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1291_
timestamp 1688980957
transform -1 0 15640 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1292_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__nand3b_2  _1293_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1294_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _1295_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15824 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__and2b_1  _1296_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14536 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1297_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16100 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1298_
timestamp 1688980957
transform 1 0 18768 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_4  _1299_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18768 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__or4bb_1  _1300_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15088 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o221ai_4  _1301_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_8  _1302_
timestamp 1688980957
transform -1 0 16468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__a221oi_2  _1303_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16928 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1304_
timestamp 1688980957
transform 1 0 20700 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1305_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1306_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21252 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1307_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20884 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1308_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20424 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1309_
timestamp 1688980957
transform 1 0 20792 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1688980957
transform -1 0 14536 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1311_
timestamp 1688980957
transform -1 0 14260 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  _1312_
timestamp 1688980957
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1313_
timestamp 1688980957
transform -1 0 18216 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1314_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17020 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1315_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12052 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1316_
timestamp 1688980957
transform 1 0 12512 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1317_
timestamp 1688980957
transform 1 0 15364 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1318_
timestamp 1688980957
transform 1 0 16100 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1319_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17296 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1320_
timestamp 1688980957
transform 1 0 16560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_4  _1321_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18308 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_1  _1322_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20240 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1323_
timestamp 1688980957
transform -1 0 20056 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _1324_
timestamp 1688980957
transform 1 0 18676 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _1325_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19504 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1326_
timestamp 1688980957
transform 1 0 18768 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1688980957
transform 1 0 17756 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1328_
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1329_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__o211a_1  _1330_
timestamp 1688980957
transform -1 0 18676 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1331_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19780 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_8  _1332_
timestamp 1688980957
transform 1 0 18216 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_4  _1333_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28796 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _1334_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15640 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_8  _1335_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__or3_4  _1336_
timestamp 1688980957
transform -1 0 14628 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1337_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15364 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_4  _1338_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14720 0 1 22848
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_1  _1339_
timestamp 1688980957
transform 1 0 12880 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1340_
timestamp 1688980957
transform 1 0 13984 0 -1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__o2bb2a_2  _1341_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1342_
timestamp 1688980957
transform 1 0 14168 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _1343_
timestamp 1688980957
transform 1 0 13524 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1344_
timestamp 1688980957
transform 1 0 15364 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__a221o_1  _1345_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27232 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1346_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28520 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1347_
timestamp 1688980957
transform -1 0 30268 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1348_
timestamp 1688980957
transform 1 0 29900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1349_
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_8  _1350_
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_2  _1351_
timestamp 1688980957
transform 1 0 16100 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1352_
timestamp 1688980957
transform -1 0 19044 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _1353_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1354_
timestamp 1688980957
transform -1 0 12328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_4  _1355_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_4  _1356_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16192 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1357_
timestamp 1688980957
transform 1 0 17296 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1358_
timestamp 1688980957
transform -1 0 20424 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1359_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19872 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _1360_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_8  _1361_
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  _1362_
timestamp 1688980957
transform 1 0 16100 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__o22ai_4  _1363_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20700 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  _1364_
timestamp 1688980957
transform 1 0 20884 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__a21oi_4  _1365_
timestamp 1688980957
transform -1 0 18124 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _1366_
timestamp 1688980957
transform -1 0 20056 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1367_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24840 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_8  _1368_
timestamp 1688980957
transform 1 0 20700 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__a211o_1  _1369_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26772 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1370_
timestamp 1688980957
transform 1 0 26036 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1371_
timestamp 1688980957
transform 1 0 25668 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1372_
timestamp 1688980957
transform -1 0 30728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1373_
timestamp 1688980957
transform -1 0 29900 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1374_
timestamp 1688980957
transform -1 0 30452 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1375_
timestamp 1688980957
transform 1 0 29624 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1376_
timestamp 1688980957
transform 1 0 30268 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1377_
timestamp 1688980957
transform -1 0 32016 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1378_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1379_
timestamp 1688980957
transform 1 0 25668 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1380_
timestamp 1688980957
transform 1 0 26220 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1381_
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1382_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 36064 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _1384_
timestamp 1688980957
transform 1 0 30360 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1385_
timestamp 1688980957
transform -1 0 32016 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1386_
timestamp 1688980957
transform -1 0 33672 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1387_
timestamp 1688980957
transform 1 0 25392 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1388_
timestamp 1688980957
transform 1 0 26036 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1389_
timestamp 1688980957
transform -1 0 26680 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1390_
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1391_
timestamp 1688980957
transform -1 0 36616 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1392_
timestamp 1688980957
transform 1 0 36616 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1393_
timestamp 1688980957
transform -1 0 37076 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1394_
timestamp 1688980957
transform 1 0 36616 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1395_
timestamp 1688980957
transform 1 0 30452 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1396_
timestamp 1688980957
transform -1 0 32016 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1397_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33672 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1398_
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1399_
timestamp 1688980957
transform -1 0 26680 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1400_
timestamp 1688980957
transform 1 0 25392 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1401_
timestamp 1688980957
transform 1 0 24840 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1402_
timestamp 1688980957
transform 1 0 25024 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1403_
timestamp 1688980957
transform -1 0 33672 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1404_
timestamp 1688980957
transform 1 0 27140 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1405_
timestamp 1688980957
transform -1 0 28980 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1406_
timestamp 1688980957
transform -1 0 30728 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1407_
timestamp 1688980957
transform -1 0 25944 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1408_
timestamp 1688980957
transform 1 0 24748 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1409_
timestamp 1688980957
transform -1 0 25300 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1410_
timestamp 1688980957
transform 1 0 25024 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1411_
timestamp 1688980957
transform 1 0 31004 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1412_
timestamp 1688980957
transform 1 0 31004 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1413_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31464 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1414_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1415_
timestamp 1688980957
transform -1 0 18584 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1416_
timestamp 1688980957
transform 1 0 17296 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _1417_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1418_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15088 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_4  _1419_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17296 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_2  _1420_
timestamp 1688980957
transform -1 0 17572 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1421_
timestamp 1688980957
transform -1 0 23460 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _1422_
timestamp 1688980957
transform 1 0 15732 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1423_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17756 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _1424_
timestamp 1688980957
transform -1 0 17112 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1425_
timestamp 1688980957
transform 1 0 20700 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1426_
timestamp 1688980957
transform 1 0 21896 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1427_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_4  _1428_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17940 0 -1 25024
box -38 -48 1326 592
use sky130_fd_sc_hd__nor4_1  _1429_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15640 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1430_
timestamp 1688980957
transform 1 0 22632 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1431_
timestamp 1688980957
transform 1 0 21344 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_2  _1432_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1433_
timestamp 1688980957
transform 1 0 11684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1435_
timestamp 1688980957
transform 1 0 12236 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1436_
timestamp 1688980957
transform 1 0 18400 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1437_
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1438_
timestamp 1688980957
transform 1 0 22080 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1439_
timestamp 1688980957
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1440_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1441_
timestamp 1688980957
transform 1 0 18308 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _1442_
timestamp 1688980957
transform -1 0 17572 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1443_
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1444_
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _1445_
timestamp 1688980957
transform 1 0 18308 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1446_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16928 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1447_
timestamp 1688980957
transform 1 0 23184 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1448_
timestamp 1688980957
transform 1 0 23736 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1449_
timestamp 1688980957
transform 1 0 17848 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1450_
timestamp 1688980957
transform 1 0 20424 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1451_
timestamp 1688980957
transform 1 0 17296 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1452_
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1453_
timestamp 1688980957
transform 1 0 23368 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1454_
timestamp 1688980957
transform 1 0 24472 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1455_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25668 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 1688980957
transform 1 0 20148 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1457_
timestamp 1688980957
transform 1 0 20976 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1458_
timestamp 1688980957
transform 1 0 20332 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1459_
timestamp 1688980957
transform 1 0 25208 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1460_
timestamp 1688980957
transform 1 0 28244 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1461_
timestamp 1688980957
transform -1 0 32384 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1462_
timestamp 1688980957
transform -1 0 32844 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1463_
timestamp 1688980957
transform 1 0 32844 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1464_
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1465_
timestamp 1688980957
transform 1 0 13524 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1466_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1467_
timestamp 1688980957
transform -1 0 15732 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1468_
timestamp 1688980957
transform -1 0 15088 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1469_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1470_
timestamp 1688980957
transform 1 0 12236 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1471_
timestamp 1688980957
transform 1 0 12420 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1472_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1473_
timestamp 1688980957
transform 1 0 17940 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _1474_
timestamp 1688980957
transform -1 0 21528 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1475_
timestamp 1688980957
transform -1 0 17296 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1476_
timestamp 1688980957
transform 1 0 16652 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1477_
timestamp 1688980957
transform 1 0 16008 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1478_
timestamp 1688980957
transform 1 0 16836 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1479_
timestamp 1688980957
transform 1 0 16100 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1480_
timestamp 1688980957
transform 1 0 17664 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1481_
timestamp 1688980957
transform -1 0 19228 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1482_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1483_
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1484_
timestamp 1688980957
transform -1 0 18124 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1485_
timestamp 1688980957
transform -1 0 18492 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_2  _1486_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18952 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1487_
timestamp 1688980957
transform -1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_4  _1488_
timestamp 1688980957
transform -1 0 19504 0 -1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _1489_
timestamp 1688980957
transform -1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1490_
timestamp 1688980957
transform -1 0 17296 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1491_
timestamp 1688980957
transform 1 0 16560 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1492_
timestamp 1688980957
transform 1 0 16100 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1493_
timestamp 1688980957
transform 1 0 17388 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1494_
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1495_
timestamp 1688980957
transform 1 0 17664 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1496_
timestamp 1688980957
transform 1 0 18492 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1497_
timestamp 1688980957
transform -1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1498_
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1499_
timestamp 1688980957
transform 1 0 18124 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1500_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18952 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1501_
timestamp 1688980957
transform -1 0 18768 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1502_
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1503_
timestamp 1688980957
transform 1 0 13064 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1504_
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1505_
timestamp 1688980957
transform -1 0 16376 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1506_
timestamp 1688980957
transform -1 0 15732 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1507_
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1508_
timestamp 1688980957
transform 1 0 11592 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1509_
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1510_
timestamp 1688980957
transform 1 0 13248 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1511_
timestamp 1688980957
transform 1 0 17572 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1512_
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1513_
timestamp 1688980957
transform 1 0 28980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1514_
timestamp 1688980957
transform 1 0 13984 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1515_
timestamp 1688980957
transform 1 0 13156 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1516_
timestamp 1688980957
transform -1 0 15180 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1517_
timestamp 1688980957
transform -1 0 20516 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1518_
timestamp 1688980957
transform 1 0 18400 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19596 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1520_
timestamp 1688980957
transform 1 0 20700 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1521_
timestamp 1688980957
transform -1 0 12236 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1522_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11592 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1523_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19964 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_4  _1524_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20700 0 -1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _1525_
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1526_
timestamp 1688980957
transform -1 0 18032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1527_
timestamp 1688980957
transform -1 0 18768 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _1528_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1529_
timestamp 1688980957
transform -1 0 17480 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1530_
timestamp 1688980957
transform 1 0 15364 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1531_
timestamp 1688980957
transform -1 0 16744 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a2111oi_1  _1532_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1533_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18676 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1534_
timestamp 1688980957
transform 1 0 17204 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1535_
timestamp 1688980957
transform 1 0 17664 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _1536_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _1537_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1538_
timestamp 1688980957
transform 1 0 18032 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1539_
timestamp 1688980957
transform 1 0 19320 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1540_
timestamp 1688980957
transform 1 0 18308 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1541_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1542_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 1688980957
transform -1 0 22816 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1544_
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1545_
timestamp 1688980957
transform 1 0 22172 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1546_
timestamp 1688980957
transform 1 0 20240 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp 1688980957
transform 1 0 20792 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1548_
timestamp 1688980957
transform -1 0 23920 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1549_
timestamp 1688980957
transform 1 0 22264 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1550_
timestamp 1688980957
transform 1 0 20424 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1551_
timestamp 1688980957
transform -1 0 21804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1552_
timestamp 1688980957
transform 1 0 20516 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1553_
timestamp 1688980957
transform -1 0 22172 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_1  _1554_
timestamp 1688980957
transform 1 0 18492 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1555_
timestamp 1688980957
transform -1 0 19872 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _1556_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1557_
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1558_
timestamp 1688980957
transform 1 0 19504 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1559_
timestamp 1688980957
transform 1 0 18676 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1560_
timestamp 1688980957
transform 1 0 18308 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1561_
timestamp 1688980957
transform -1 0 13524 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1562_
timestamp 1688980957
transform 1 0 12144 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1563_
timestamp 1688980957
transform 1 0 12788 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1564_
timestamp 1688980957
transform 1 0 18216 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1565_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19320 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1566_
timestamp 1688980957
transform 1 0 19504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1567_
timestamp 1688980957
transform -1 0 20056 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1568_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1569_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20700 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1570_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1571_
timestamp 1688980957
transform -1 0 23736 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1572_
timestamp 1688980957
transform 1 0 20608 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1573_
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1574_
timestamp 1688980957
transform -1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1575_
timestamp 1688980957
transform -1 0 23276 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1576_
timestamp 1688980957
transform 1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1577_
timestamp 1688980957
transform 1 0 20700 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _1578_
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_2  _1579_
timestamp 1688980957
transform 1 0 26404 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1580_
timestamp 1688980957
transform -1 0 24380 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1581_
timestamp 1688980957
transform -1 0 25024 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp 1688980957
transform 1 0 23460 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1583_
timestamp 1688980957
transform 1 0 22724 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1584_
timestamp 1688980957
transform 1 0 23184 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1585_
timestamp 1688980957
transform -1 0 24564 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1586_
timestamp 1688980957
transform 1 0 23368 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1587_
timestamp 1688980957
transform 1 0 19044 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1588_
timestamp 1688980957
transform -1 0 20148 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1589_
timestamp 1688980957
transform 1 0 20148 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1590_
timestamp 1688980957
transform -1 0 20148 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1591_
timestamp 1688980957
transform 1 0 22816 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1592_
timestamp 1688980957
transform 1 0 28704 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1593_
timestamp 1688980957
transform 1 0 28796 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1594_
timestamp 1688980957
transform 1 0 31832 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1595_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30268 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1596_
timestamp 1688980957
transform -1 0 24196 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1597_
timestamp 1688980957
transform 1 0 20792 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1598_
timestamp 1688980957
transform 1 0 21896 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1599_
timestamp 1688980957
transform 1 0 22816 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1600_
timestamp 1688980957
transform -1 0 24012 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1601_
timestamp 1688980957
transform 1 0 23184 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1602_
timestamp 1688980957
transform 1 0 23368 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1603_
timestamp 1688980957
transform -1 0 24196 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1604_
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1605_
timestamp 1688980957
transform -1 0 24840 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1606_
timestamp 1688980957
transform 1 0 23644 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 1688980957
transform 1 0 23276 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1608_
timestamp 1688980957
transform 1 0 24012 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1609_
timestamp 1688980957
transform 1 0 23368 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1610_
timestamp 1688980957
transform 1 0 23552 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1611_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24472 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1612_
timestamp 1688980957
transform 1 0 23552 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1613_
timestamp 1688980957
transform 1 0 20976 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1614_
timestamp 1688980957
transform 1 0 21896 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1615_
timestamp 1688980957
transform -1 0 23184 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _1616_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24012 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _1617_
timestamp 1688980957
transform 1 0 24104 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__a22oi_1  _1618_
timestamp 1688980957
transform -1 0 14812 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1619_
timestamp 1688980957
transform 1 0 13340 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1620_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1621_
timestamp 1688980957
transform 1 0 15272 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1622_
timestamp 1688980957
transform 1 0 13248 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1623_
timestamp 1688980957
transform 1 0 13524 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1624_
timestamp 1688980957
transform -1 0 13432 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1688980957
transform 1 0 11224 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_2  _1626_
timestamp 1688980957
transform 1 0 11868 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _1627_
timestamp 1688980957
transform 1 0 26128 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1628_
timestamp 1688980957
transform -1 0 19136 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1629_
timestamp 1688980957
transform -1 0 18768 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1630_
timestamp 1688980957
transform 1 0 15916 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1631_
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1632_
timestamp 1688980957
transform 1 0 17204 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1633_
timestamp 1688980957
transform 1 0 17480 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1634_
timestamp 1688980957
transform 1 0 17756 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1635_
timestamp 1688980957
transform 1 0 18308 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1636_
timestamp 1688980957
transform 1 0 15916 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1637_
timestamp 1688980957
transform 1 0 16744 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1638_
timestamp 1688980957
transform 1 0 18216 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_4  _1639_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19136 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_2  _1640_
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1641_
timestamp 1688980957
transform -1 0 30636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1642_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31372 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1643_
timestamp 1688980957
transform 1 0 25944 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1644_
timestamp 1688980957
transform 1 0 26036 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1645_
timestamp 1688980957
transform -1 0 27600 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1646_
timestamp 1688980957
transform 1 0 30176 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1647_
timestamp 1688980957
transform -1 0 30636 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1648_
timestamp 1688980957
transform -1 0 33212 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1649_
timestamp 1688980957
transform 1 0 31188 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1650_
timestamp 1688980957
transform -1 0 31648 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1651_
timestamp 1688980957
transform -1 0 33028 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1652_
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1653_
timestamp 1688980957
transform 1 0 36064 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1654_
timestamp 1688980957
transform 1 0 35420 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1655_
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1656_
timestamp 1688980957
transform 1 0 36156 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1657_
timestamp 1688980957
transform 1 0 35144 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1658_
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1659_
timestamp 1688980957
transform -1 0 32016 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1660_
timestamp 1688980957
transform -1 0 32844 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1688980957
transform -1 0 26588 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1662_
timestamp 1688980957
transform -1 0 26680 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1663_
timestamp 1688980957
transform -1 0 27692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1664_
timestamp 1688980957
transform 1 0 27692 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1665_
timestamp 1688980957
transform 1 0 33028 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1666_
timestamp 1688980957
transform 1 0 33580 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1667_
timestamp 1688980957
transform -1 0 34132 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1668_
timestamp 1688980957
transform 1 0 34132 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1669_
timestamp 1688980957
transform 1 0 30360 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1670_
timestamp 1688980957
transform 1 0 31096 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_2  _1671_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31096 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1672_
timestamp 1688980957
transform -1 0 26404 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1673_
timestamp 1688980957
transform -1 0 26128 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1674_
timestamp 1688980957
transform -1 0 26864 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1675_
timestamp 1688980957
transform 1 0 27048 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1676_
timestamp 1688980957
transform -1 0 31648 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1677_
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1678_
timestamp 1688980957
transform 1 0 32200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1679_
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1680_
timestamp 1688980957
transform -1 0 33580 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1681_
timestamp 1688980957
transform 1 0 32568 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1682_
timestamp 1688980957
transform 1 0 32200 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1683_
timestamp 1688980957
transform -1 0 31004 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1684_
timestamp 1688980957
transform 1 0 29624 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1685_
timestamp 1688980957
transform 1 0 30360 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1686_
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1687_
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1688_
timestamp 1688980957
transform 1 0 25484 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1689_
timestamp 1688980957
transform -1 0 26036 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1690_
timestamp 1688980957
transform 1 0 25760 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1691_
timestamp 1688980957
transform 1 0 28980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1692_
timestamp 1688980957
transform 1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1688980957
transform 1 0 29716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1694_
timestamp 1688980957
transform 1 0 29992 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1695_
timestamp 1688980957
transform 1 0 30176 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1696_
timestamp 1688980957
transform 1 0 20332 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1697_
timestamp 1688980957
transform 1 0 19596 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1698_
timestamp 1688980957
transform 1 0 20332 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1699_
timestamp 1688980957
transform 1 0 20240 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1700_
timestamp 1688980957
transform 1 0 20976 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__and3b_2  _1701_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1702_
timestamp 1688980957
transform -1 0 20608 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1703_
timestamp 1688980957
transform 1 0 19688 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1704_
timestamp 1688980957
transform 1 0 19688 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__o211ai_4  _1705_
timestamp 1688980957
transform 1 0 20148 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_8  _1706_
timestamp 1688980957
transform -1 0 23276 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_2  _1707_
timestamp 1688980957
transform 1 0 27876 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1708_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30176 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1709_
timestamp 1688980957
transform 1 0 35144 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1710_
timestamp 1688980957
transform 1 0 33856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1711_
timestamp 1688980957
transform 1 0 34684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1712_
timestamp 1688980957
transform 1 0 32016 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1713_
timestamp 1688980957
transform -1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1714_
timestamp 1688980957
transform 1 0 21160 0 1 4352
box -38 -48 2062 592
use sky130_fd_sc_hd__o211a_1  _1715_
timestamp 1688980957
transform -1 0 18860 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1716_
timestamp 1688980957
transform 1 0 20240 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1717_
timestamp 1688980957
transform -1 0 21712 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1718_
timestamp 1688980957
transform 1 0 26404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1719_
timestamp 1688980957
transform 1 0 25576 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1720_
timestamp 1688980957
transform -1 0 26680 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1721_
timestamp 1688980957
transform -1 0 29440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1722_
timestamp 1688980957
transform -1 0 29900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1723_
timestamp 1688980957
transform 1 0 25208 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1724_
timestamp 1688980957
transform 1 0 25484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1725_
timestamp 1688980957
transform 1 0 25208 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1726_
timestamp 1688980957
transform 1 0 26404 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1727_
timestamp 1688980957
transform -1 0 27324 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1728_
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _1729_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22908 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1730_
timestamp 1688980957
transform -1 0 27968 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1731_
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1732_
timestamp 1688980957
transform -1 0 26036 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1733_
timestamp 1688980957
transform -1 0 26864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1734_
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1735_
timestamp 1688980957
transform -1 0 25944 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1736_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29256 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1737_
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1738_
timestamp 1688980957
transform 1 0 33304 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1739_
timestamp 1688980957
transform -1 0 34684 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1740_
timestamp 1688980957
transform 1 0 34960 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1741_
timestamp 1688980957
transform -1 0 36156 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1742_
timestamp 1688980957
transform 1 0 35512 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1743_
timestamp 1688980957
transform 1 0 31648 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1744_
timestamp 1688980957
transform -1 0 33580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1745_
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1746_
timestamp 1688980957
transform 1 0 29716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1747_
timestamp 1688980957
transform 1 0 29532 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1748_
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _1749_
timestamp 1688980957
transform 1 0 22540 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1750_
timestamp 1688980957
transform 1 0 30084 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_4  _1751_
timestamp 1688980957
transform 1 0 30268 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1752_
timestamp 1688980957
transform 1 0 29072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1753_
timestamp 1688980957
transform 1 0 30544 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1754_
timestamp 1688980957
transform 1 0 31004 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1755_
timestamp 1688980957
transform 1 0 31464 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1756_
timestamp 1688980957
transform 1 0 29348 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1757_
timestamp 1688980957
transform 1 0 29900 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1758_
timestamp 1688980957
transform -1 0 33028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1759_
timestamp 1688980957
transform -1 0 33672 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1760_
timestamp 1688980957
transform -1 0 33304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1761_
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1762_
timestamp 1688980957
transform 1 0 31648 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1763_
timestamp 1688980957
transform 1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1764_
timestamp 1688980957
transform 1 0 19780 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1765_
timestamp 1688980957
transform 1 0 19504 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1766_
timestamp 1688980957
transform -1 0 20332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1767_
timestamp 1688980957
transform 1 0 19596 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1768_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19964 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1769_
timestamp 1688980957
transform -1 0 25576 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1770_
timestamp 1688980957
transform -1 0 28980 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1771_
timestamp 1688980957
transform -1 0 27140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1772_
timestamp 1688980957
transform 1 0 30912 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1773_
timestamp 1688980957
transform 1 0 32108 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1774_
timestamp 1688980957
transform -1 0 33396 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1775_
timestamp 1688980957
transform -1 0 32844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1776_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33580 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1777_
timestamp 1688980957
transform -1 0 34132 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1778_
timestamp 1688980957
transform -1 0 33488 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _1779_
timestamp 1688980957
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1780_
timestamp 1688980957
transform -1 0 21436 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1781_
timestamp 1688980957
transform -1 0 29072 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1782_
timestamp 1688980957
transform -1 0 32568 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1783_
timestamp 1688980957
transform -1 0 33028 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1784_
timestamp 1688980957
transform 1 0 28888 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1785_
timestamp 1688980957
transform 1 0 28888 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1786_
timestamp 1688980957
transform -1 0 29348 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1787_
timestamp 1688980957
transform -1 0 29072 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1788_
timestamp 1688980957
transform 1 0 30452 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1789_
timestamp 1688980957
transform 1 0 32568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1790_
timestamp 1688980957
transform -1 0 30176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1791_
timestamp 1688980957
transform -1 0 32752 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1792_
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1793_
timestamp 1688980957
transform 1 0 29992 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1794_
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1795_
timestamp 1688980957
transform 1 0 18952 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1796_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1797_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1798_
timestamp 1688980957
transform 1 0 20792 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1799_
timestamp 1688980957
transform 1 0 21528 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1800_
timestamp 1688980957
transform 1 0 22172 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1801_
timestamp 1688980957
transform 1 0 25576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1802_
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1803_
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1804_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 31924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1805_
timestamp 1688980957
transform -1 0 31464 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1806_
timestamp 1688980957
transform -1 0 29808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1807_
timestamp 1688980957
transform -1 0 21528 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _1808_
timestamp 1688980957
transform 1 0 22172 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a2111oi_1  _1809_
timestamp 1688980957
transform 1 0 28060 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1810_
timestamp 1688980957
transform -1 0 28796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1811_
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1812_
timestamp 1688980957
transform 1 0 32108 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1813_
timestamp 1688980957
transform -1 0 30912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1814_
timestamp 1688980957
transform 1 0 27968 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1815_
timestamp 1688980957
transform -1 0 27876 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1816_
timestamp 1688980957
transform 1 0 20424 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1817_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21896 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1818_
timestamp 1688980957
transform -1 0 23828 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1819_
timestamp 1688980957
transform 1 0 22448 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1820_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20608 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1821_
timestamp 1688980957
transform -1 0 23276 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1822_
timestamp 1688980957
transform 1 0 22356 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1823_
timestamp 1688980957
transform 1 0 33028 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1824_
timestamp 1688980957
transform -1 0 23552 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_4  _1825_
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1826_
timestamp 1688980957
transform 1 0 26312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1827_
timestamp 1688980957
transform 1 0 25392 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1828_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1829_
timestamp 1688980957
transform -1 0 21804 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1830_
timestamp 1688980957
transform 1 0 19504 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1831_
timestamp 1688980957
transform 1 0 24840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1832_
timestamp 1688980957
transform 1 0 23460 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1833_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25208 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1834_
timestamp 1688980957
transform 1 0 24932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1835_
timestamp 1688980957
transform -1 0 24932 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1836_
timestamp 1688980957
transform -1 0 25392 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1837_
timestamp 1688980957
transform -1 0 27508 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1838_
timestamp 1688980957
transform -1 0 29348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1839_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27508 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1840_
timestamp 1688980957
transform -1 0 25024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1841_
timestamp 1688980957
transform 1 0 25668 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1842_
timestamp 1688980957
transform -1 0 19596 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1843_
timestamp 1688980957
transform -1 0 20608 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1844_
timestamp 1688980957
transform 1 0 20148 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _1845_
timestamp 1688980957
transform 1 0 20608 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1846_
timestamp 1688980957
transform -1 0 19964 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1847_
timestamp 1688980957
transform -1 0 20240 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1848_
timestamp 1688980957
transform 1 0 20516 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1849_
timestamp 1688980957
transform 1 0 22264 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _1850_
timestamp 1688980957
transform 1 0 21344 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1851_
timestamp 1688980957
transform -1 0 14812 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1852_
timestamp 1688980957
transform -1 0 16560 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1853_
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1854_
timestamp 1688980957
transform 1 0 16744 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1855_
timestamp 1688980957
transform -1 0 16376 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1856_
timestamp 1688980957
transform 1 0 15456 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1857_
timestamp 1688980957
transform 1 0 14168 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1858_
timestamp 1688980957
transform 1 0 14812 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_4  _1859_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22908 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_4  _1860_
timestamp 1688980957
transform -1 0 25576 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1861_
timestamp 1688980957
transform -1 0 33856 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1862_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 34132 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1863_
timestamp 1688980957
transform -1 0 33212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1864_
timestamp 1688980957
transform -1 0 33212 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1865_
timestamp 1688980957
transform 1 0 28152 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1866_
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1867_
timestamp 1688980957
transform 1 0 31464 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1868_
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1869_
timestamp 1688980957
transform 1 0 30176 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1870_
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _1871_
timestamp 1688980957
transform 1 0 23552 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _1872_
timestamp 1688980957
transform 1 0 23276 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1873_
timestamp 1688980957
transform 1 0 26036 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1874_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25944 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1875_
timestamp 1688980957
transform -1 0 26956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1876_
timestamp 1688980957
transform -1 0 27508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1877_
timestamp 1688980957
transform 1 0 30176 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1878_
timestamp 1688980957
transform -1 0 32016 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1879_
timestamp 1688980957
transform -1 0 31464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1880_
timestamp 1688980957
transform 1 0 30728 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_2  _1881_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30728 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1882_
timestamp 1688980957
transform -1 0 27876 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1883_
timestamp 1688980957
transform -1 0 27416 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1884_
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1885_
timestamp 1688980957
transform -1 0 26864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1886_
timestamp 1688980957
transform 1 0 31464 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1887_
timestamp 1688980957
transform 1 0 31096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1888_
timestamp 1688980957
transform 1 0 32384 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1889_
timestamp 1688980957
transform 1 0 25392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1890_
timestamp 1688980957
transform 1 0 26864 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1891_
timestamp 1688980957
transform -1 0 26864 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1892_
timestamp 1688980957
transform -1 0 27692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1893_
timestamp 1688980957
transform 1 0 30084 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1894_
timestamp 1688980957
transform 1 0 32844 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1895_
timestamp 1688980957
transform -1 0 28704 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1896_
timestamp 1688980957
transform -1 0 33028 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1897_
timestamp 1688980957
transform 1 0 32384 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1898_
timestamp 1688980957
transform -1 0 32016 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1899_
timestamp 1688980957
transform 1 0 33120 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1900_
timestamp 1688980957
transform -1 0 33764 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1901_
timestamp 1688980957
transform -1 0 32384 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1902_
timestamp 1688980957
transform 1 0 32292 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1903_
timestamp 1688980957
transform -1 0 32200 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1904_
timestamp 1688980957
transform 1 0 32476 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1905_
timestamp 1688980957
transform 1 0 32476 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1906_
timestamp 1688980957
transform 1 0 27968 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1907_
timestamp 1688980957
transform 1 0 30084 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1908_
timestamp 1688980957
transform -1 0 29900 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1909_
timestamp 1688980957
transform 1 0 30912 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1910_
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1911_
timestamp 1688980957
transform -1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1912_
timestamp 1688980957
transform 1 0 30084 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1913_
timestamp 1688980957
transform 1 0 23828 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1914_
timestamp 1688980957
transform -1 0 23828 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1915_
timestamp 1688980957
transform 1 0 21528 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1916_
timestamp 1688980957
transform -1 0 24380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1917_
timestamp 1688980957
transform 1 0 25944 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1918_
timestamp 1688980957
transform 1 0 27600 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1919_
timestamp 1688980957
transform 1 0 26772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1920_
timestamp 1688980957
transform 1 0 24380 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1921_
timestamp 1688980957
transform -1 0 27692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1922_
timestamp 1688980957
transform -1 0 28888 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_2  _1923_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__o211a_1  _1924_
timestamp 1688980957
transform 1 0 31464 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1925_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30728 0 -1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _1926_
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1927_
timestamp 1688980957
transform -1 0 34040 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1928_
timestamp 1688980957
transform 1 0 33028 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1929_
timestamp 1688980957
transform 1 0 28612 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1930_
timestamp 1688980957
transform 1 0 34224 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1931_
timestamp 1688980957
transform -1 0 34592 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1932_
timestamp 1688980957
transform 1 0 26128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1933_
timestamp 1688980957
transform 1 0 27140 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1934_
timestamp 1688980957
transform -1 0 27968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1935_
timestamp 1688980957
transform -1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1936_
timestamp 1688980957
transform -1 0 28060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1937_
timestamp 1688980957
transform 1 0 27600 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_1  _1938_
timestamp 1688980957
transform -1 0 25852 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1939_
timestamp 1688980957
transform -1 0 26588 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1940_
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1941_
timestamp 1688980957
transform 1 0 26956 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1942_
timestamp 1688980957
transform 1 0 27508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1943_
timestamp 1688980957
transform -1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1944_
timestamp 1688980957
transform 1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1945_
timestamp 1688980957
transform -1 0 28888 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1946_
timestamp 1688980957
transform -1 0 36800 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1947_
timestamp 1688980957
transform 1 0 35420 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1948_
timestamp 1688980957
transform -1 0 35696 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _1949_
timestamp 1688980957
transform -1 0 35420 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1950_
timestamp 1688980957
transform 1 0 27232 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1951_
timestamp 1688980957
transform -1 0 34592 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1952_
timestamp 1688980957
transform -1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1953_
timestamp 1688980957
transform 1 0 22356 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1954_
timestamp 1688980957
transform 1 0 23000 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1955_
timestamp 1688980957
transform -1 0 23552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1956_
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1957_
timestamp 1688980957
transform 1 0 19964 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1958_
timestamp 1688980957
transform 1 0 20884 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1959_
timestamp 1688980957
transform 1 0 25392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1960_
timestamp 1688980957
transform -1 0 19044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1961_
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1962_
timestamp 1688980957
transform 1 0 25392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1963_
timestamp 1688980957
transform -1 0 25392 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1964_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1965_
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1966_
timestamp 1688980957
transform 1 0 23368 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_4  _1967_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23920 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1968_
timestamp 1688980957
transform 1 0 35788 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1969_
timestamp 1688980957
transform 1 0 35512 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1970_
timestamp 1688980957
transform 1 0 36340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1971_
timestamp 1688980957
transform 1 0 34776 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1972_
timestamp 1688980957
transform -1 0 25760 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1973_
timestamp 1688980957
transform 1 0 24840 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1974_
timestamp 1688980957
transform -1 0 34868 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1975_
timestamp 1688980957
transform -1 0 34960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1976_
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1977_
timestamp 1688980957
transform 1 0 21896 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1978_
timestamp 1688980957
transform 1 0 19688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1979_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1980_
timestamp 1688980957
transform -1 0 22448 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1981_
timestamp 1688980957
transform 1 0 19688 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1982_
timestamp 1688980957
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1983_
timestamp 1688980957
transform -1 0 22908 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1984_
timestamp 1688980957
transform 1 0 22908 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1985_
timestamp 1688980957
transform 1 0 23000 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1986_
timestamp 1688980957
transform 1 0 21804 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1987_
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_4  _1988_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__a21oi_1  _1989_
timestamp 1688980957
transform -1 0 33212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1990_
timestamp 1688980957
transform -1 0 34776 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1991_
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1992_
timestamp 1688980957
transform -1 0 35420 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1993_
timestamp 1688980957
transform -1 0 33764 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1994_
timestamp 1688980957
transform 1 0 27232 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1995_
timestamp 1688980957
transform -1 0 34684 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1996_
timestamp 1688980957
transform -1 0 34960 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1997_
timestamp 1688980957
transform -1 0 21712 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1998_
timestamp 1688980957
transform -1 0 20884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1999_
timestamp 1688980957
transform -1 0 20516 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2000_
timestamp 1688980957
transform 1 0 21620 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _2001_
timestamp 1688980957
transform 1 0 20884 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2002_
timestamp 1688980957
transform 1 0 22724 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2003_
timestamp 1688980957
transform 1 0 22448 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2004_
timestamp 1688980957
transform 1 0 21988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2005_
timestamp 1688980957
transform 1 0 24564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2006_
timestamp 1688980957
transform 1 0 21344 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2007_
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _2008_
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2009_
timestamp 1688980957
transform -1 0 30544 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2010_
timestamp 1688980957
transform -1 0 32568 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2011_
timestamp 1688980957
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2012_
timestamp 1688980957
transform -1 0 32844 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _2013_
timestamp 1688980957
transform 1 0 32844 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2014_
timestamp 1688980957
transform -1 0 27048 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2015_
timestamp 1688980957
transform -1 0 29164 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2016_
timestamp 1688980957
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2017_
timestamp 1688980957
transform 1 0 23092 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2018_
timestamp 1688980957
transform 1 0 27600 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2019_
timestamp 1688980957
transform 1 0 29164 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2020_
timestamp 1688980957
transform -1 0 29072 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2021_
timestamp 1688980957
transform 1 0 27324 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2022_
timestamp 1688980957
transform -1 0 26864 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2023_
timestamp 1688980957
transform 1 0 28060 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2024_
timestamp 1688980957
transform 1 0 28060 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2025_
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2026_
timestamp 1688980957
transform -1 0 29348 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2027_
timestamp 1688980957
transform -1 0 28336 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2028_
timestamp 1688980957
transform 1 0 28336 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2029_
timestamp 1688980957
transform -1 0 30360 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2030_
timestamp 1688980957
transform 1 0 29808 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2031_
timestamp 1688980957
transform 1 0 28428 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2032_
timestamp 1688980957
transform -1 0 28152 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2033_
timestamp 1688980957
transform 1 0 27784 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2034_
timestamp 1688980957
transform 1 0 27968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2035_
timestamp 1688980957
transform -1 0 13984 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _2036_
timestamp 1688980957
transform -1 0 14904 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and4_2  _2037_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _2038_
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2039_
timestamp 1688980957
transform 1 0 24288 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2040_
timestamp 1688980957
transform -1 0 23092 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2041_
timestamp 1688980957
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2042_
timestamp 1688980957
transform -1 0 22632 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _2043_
timestamp 1688980957
transform 1 0 22172 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_4  _2044_
timestamp 1688980957
transform 1 0 22632 0 -1 23936
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2045_
timestamp 1688980957
transform 1 0 19412 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2046_
timestamp 1688980957
transform -1 0 19688 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2047_
timestamp 1688980957
transform 1 0 9568 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2048_
timestamp 1688980957
transform 1 0 10212 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2049_
timestamp 1688980957
transform 1 0 9752 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2050_
timestamp 1688980957
transform -1 0 9752 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2051_
timestamp 1688980957
transform -1 0 10212 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2052_
timestamp 1688980957
transform 1 0 9660 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2053_
timestamp 1688980957
transform -1 0 10396 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2054_
timestamp 1688980957
transform 1 0 8740 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2055_
timestamp 1688980957
transform -1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2056_
timestamp 1688980957
transform 1 0 9200 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2057_
timestamp 1688980957
transform 1 0 10120 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2058_
timestamp 1688980957
transform 1 0 9844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2059_
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2060_
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2061_
timestamp 1688980957
transform 1 0 10580 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2062_
timestamp 1688980957
transform 1 0 8740 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2063_
timestamp 1688980957
transform 1 0 9476 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2064_
timestamp 1688980957
transform 1 0 9568 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2065_
timestamp 1688980957
transform 1 0 9844 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2066_
timestamp 1688980957
transform 1 0 11960 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2067_
timestamp 1688980957
transform 1 0 10580 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2068_
timestamp 1688980957
transform -1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _2069_
timestamp 1688980957
transform -1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2070_
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _2071_
timestamp 1688980957
transform -1 0 25392 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2072_
timestamp 1688980957
transform -1 0 31372 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2073_
timestamp 1688980957
transform 1 0 31004 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2074_
timestamp 1688980957
transform 1 0 26036 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2075_
timestamp 1688980957
transform 1 0 26220 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2076_
timestamp 1688980957
transform -1 0 28980 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2077_
timestamp 1688980957
transform 1 0 28980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2078_
timestamp 1688980957
transform -1 0 33028 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2079_
timestamp 1688980957
transform 1 0 32844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2080_
timestamp 1688980957
transform -1 0 33856 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2081_
timestamp 1688980957
transform -1 0 34132 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2082_
timestamp 1688980957
transform 1 0 33212 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2083_
timestamp 1688980957
transform -1 0 33396 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2084_
timestamp 1688980957
transform -1 0 33764 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2085_
timestamp 1688980957
transform 1 0 33304 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2086_
timestamp 1688980957
transform -1 0 26864 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2087_
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2088_
timestamp 1688980957
transform 1 0 23276 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2089_
timestamp 1688980957
transform 1 0 21988 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2090_
timestamp 1688980957
transform -1 0 21528 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2091_
timestamp 1688980957
transform -1 0 12328 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2092_
timestamp 1688980957
transform -1 0 12328 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2093_
timestamp 1688980957
transform 1 0 5428 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2094_
timestamp 1688980957
transform 1 0 5428 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2095_
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2096_
timestamp 1688980957
transform 1 0 4600 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2097_
timestamp 1688980957
transform 1 0 7820 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2098_
timestamp 1688980957
transform 1 0 6440 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2099_
timestamp 1688980957
transform 1 0 11592 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2100_
timestamp 1688980957
transform 1 0 10212 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2101_
timestamp 1688980957
transform 1 0 7268 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2102_
timestamp 1688980957
transform 1 0 6532 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2103_
timestamp 1688980957
transform 1 0 9292 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2104_
timestamp 1688980957
transform 1 0 9016 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2105_
timestamp 1688980957
transform -1 0 24288 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _2106_
timestamp 1688980957
transform 1 0 23092 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2107_
timestamp 1688980957
transform 1 0 32568 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2108_
timestamp 1688980957
transform -1 0 32292 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2109_
timestamp 1688980957
transform -1 0 28152 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2110_
timestamp 1688980957
transform 1 0 28152 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2111_
timestamp 1688980957
transform -1 0 31280 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2112_
timestamp 1688980957
transform -1 0 31188 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2113_
timestamp 1688980957
transform -1 0 34592 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2114_
timestamp 1688980957
transform -1 0 34500 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2115_
timestamp 1688980957
transform -1 0 35512 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2116_
timestamp 1688980957
transform 1 0 35236 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2117_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2118_
timestamp 1688980957
transform 1 0 31464 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2119_
timestamp 1688980957
transform 1 0 31188 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2120_
timestamp 1688980957
transform 1 0 31188 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2121_
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2122_
timestamp 1688980957
transform 1 0 25944 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _2123_
timestamp 1688980957
transform -1 0 23092 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _2124_
timestamp 1688980957
transform 1 0 22356 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2125_
timestamp 1688980957
transform 1 0 20884 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2126_
timestamp 1688980957
transform 1 0 9292 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2127_
timestamp 1688980957
transform -1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2128_
timestamp 1688980957
transform 1 0 6256 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2129_
timestamp 1688980957
transform 1 0 4968 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2130_
timestamp 1688980957
transform 1 0 5428 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2131_
timestamp 1688980957
transform 1 0 4508 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2132_
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2133_
timestamp 1688980957
transform 1 0 8280 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2134_
timestamp 1688980957
transform 1 0 9568 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2135_
timestamp 1688980957
transform 1 0 8280 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2136_
timestamp 1688980957
transform 1 0 7912 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2137_
timestamp 1688980957
transform 1 0 7636 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2138_
timestamp 1688980957
transform 1 0 9200 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2139_
timestamp 1688980957
transform 1 0 7912 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2140_
timestamp 1688980957
transform -1 0 24656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2141_
timestamp 1688980957
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2142_
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2143_
timestamp 1688980957
transform 1 0 18308 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2144_
timestamp 1688980957
transform -1 0 18308 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2145_
timestamp 1688980957
transform 1 0 17664 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2146_
timestamp 1688980957
transform 1 0 17480 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _2147_
timestamp 1688980957
transform 1 0 15272 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_4  _2148_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__a31o_2  _2149_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2150_
timestamp 1688980957
transform 1 0 6900 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2151_
timestamp 1688980957
transform 1 0 5428 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2152_
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2153_
timestamp 1688980957
transform -1 0 25392 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2154_
timestamp 1688980957
transform 1 0 24104 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2155_
timestamp 1688980957
transform 1 0 23828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2156_
timestamp 1688980957
transform 1 0 22172 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2157_
timestamp 1688980957
transform 1 0 22816 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _2158_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24012 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2159_
timestamp 1688980957
transform -1 0 10488 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2160_
timestamp 1688980957
transform 1 0 9476 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2161_
timestamp 1688980957
transform -1 0 9936 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2162_
timestamp 1688980957
transform -1 0 7912 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2163_
timestamp 1688980957
transform -1 0 7360 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2164_
timestamp 1688980957
transform -1 0 8096 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2165_
timestamp 1688980957
transform 1 0 31740 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2166_
timestamp 1688980957
transform 1 0 29440 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2167_
timestamp 1688980957
transform -1 0 30360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2168_
timestamp 1688980957
transform 1 0 29992 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2169_
timestamp 1688980957
transform 1 0 23184 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2170_
timestamp 1688980957
transform 1 0 24104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2171_
timestamp 1688980957
transform 1 0 23828 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2172_
timestamp 1688980957
transform 1 0 24104 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2173_
timestamp 1688980957
transform 1 0 24748 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2174_
timestamp 1688980957
transform 1 0 33028 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2175_
timestamp 1688980957
transform 1 0 33488 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2176_
timestamp 1688980957
transform 1 0 33488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2177_
timestamp 1688980957
transform -1 0 24656 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2178_
timestamp 1688980957
transform 1 0 33856 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2179_
timestamp 1688980957
transform 1 0 34500 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2180_
timestamp 1688980957
transform -1 0 35972 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2181_
timestamp 1688980957
transform 1 0 32936 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2182_
timestamp 1688980957
transform -1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2183_
timestamp 1688980957
transform 1 0 33764 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2184_
timestamp 1688980957
transform 1 0 34408 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2185_
timestamp 1688980957
transform 1 0 34868 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2186_
timestamp 1688980957
transform 1 0 28244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2187_
timestamp 1688980957
transform 1 0 30912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2188_
timestamp 1688980957
transform 1 0 31188 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2189_
timestamp 1688980957
transform 1 0 32844 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2190_
timestamp 1688980957
transform 1 0 33764 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2191_
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2192_
timestamp 1688980957
transform -1 0 35236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2193_
timestamp 1688980957
transform 1 0 34960 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2194_
timestamp 1688980957
transform 1 0 35420 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2195_
timestamp 1688980957
transform -1 0 34592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_4  _2196_
timestamp 1688980957
transform 1 0 28152 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_1  _2197_
timestamp 1688980957
transform -1 0 28336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2198_
timestamp 1688980957
transform -1 0 28796 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2199_
timestamp 1688980957
transform 1 0 22172 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2200_
timestamp 1688980957
transform 1 0 23368 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2201_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2202_
timestamp 1688980957
transform 1 0 25024 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2203_
timestamp 1688980957
transform 1 0 25668 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2204_
timestamp 1688980957
transform 1 0 26036 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2205_
timestamp 1688980957
transform 1 0 26864 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2206_
timestamp 1688980957
transform 1 0 27968 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_4  _2207_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29256 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _2208_
timestamp 1688980957
transform 1 0 9384 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2209_
timestamp 1688980957
transform 1 0 8004 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2210_
timestamp 1688980957
transform 1 0 7728 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2211_
timestamp 1688980957
transform -1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2212_
timestamp 1688980957
transform 1 0 7636 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2213_
timestamp 1688980957
transform 1 0 30452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2214_
timestamp 1688980957
transform -1 0 30268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2215_
timestamp 1688980957
transform 1 0 29072 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2216_
timestamp 1688980957
transform 1 0 23460 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2217_
timestamp 1688980957
transform -1 0 23460 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2218_
timestamp 1688980957
transform -1 0 24564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _2219_
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _2220_
timestamp 1688980957
transform -1 0 30268 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2221_
timestamp 1688980957
transform -1 0 28980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2222_
timestamp 1688980957
transform 1 0 28428 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2223_
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _2224_
timestamp 1688980957
transform -1 0 29716 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _2225_
timestamp 1688980957
transform 1 0 28980 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2226_
timestamp 1688980957
transform -1 0 12236 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2227_
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2228_
timestamp 1688980957
transform 1 0 11040 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2229_
timestamp 1688980957
transform 1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2230_
timestamp 1688980957
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _2231_
timestamp 1688980957
transform -1 0 12972 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2232_
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2233_
timestamp 1688980957
transform -1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2234_
timestamp 1688980957
transform -1 0 15088 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _2235_
timestamp 1688980957
transform -1 0 16928 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_2  _2236_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _2237_
timestamp 1688980957
transform -1 0 14628 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2238_
timestamp 1688980957
transform 1 0 9016 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2239_
timestamp 1688980957
transform -1 0 10120 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2240_
timestamp 1688980957
transform 1 0 9384 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2241_
timestamp 1688980957
transform -1 0 10304 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _2242_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13248 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _2243_
timestamp 1688980957
transform -1 0 13616 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2244_
timestamp 1688980957
transform 1 0 8464 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2245_
timestamp 1688980957
transform 1 0 8372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2246_
timestamp 1688980957
transform -1 0 8832 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2247_
timestamp 1688980957
transform 1 0 8924 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2248_
timestamp 1688980957
transform -1 0 9660 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2249_
timestamp 1688980957
transform -1 0 9108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2250_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2251_
timestamp 1688980957
transform 1 0 7912 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2252_
timestamp 1688980957
transform -1 0 8740 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2253_
timestamp 1688980957
transform -1 0 8648 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2254_
timestamp 1688980957
transform -1 0 10396 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2255_
timestamp 1688980957
transform -1 0 8004 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2256_
timestamp 1688980957
transform -1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_2  _2257_
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _2258_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _2259_
timestamp 1688980957
transform 1 0 7452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2260_
timestamp 1688980957
transform -1 0 10212 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2261_
timestamp 1688980957
transform 1 0 8280 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _2262_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2263_
timestamp 1688980957
transform -1 0 9568 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2264_
timestamp 1688980957
transform -1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2265_
timestamp 1688980957
transform 1 0 10120 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2266_
timestamp 1688980957
transform -1 0 14352 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2267_
timestamp 1688980957
transform -1 0 14628 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _2268_
timestamp 1688980957
transform 1 0 14352 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  _2269_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7728 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2270_
timestamp 1688980957
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2271_
timestamp 1688980957
transform 1 0 15548 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2272_
timestamp 1688980957
transform 1 0 15364 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2273_
timestamp 1688980957
transform 1 0 16008 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  _2274_
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2275_
timestamp 1688980957
transform -1 0 15548 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2276_
timestamp 1688980957
transform 1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2277_
timestamp 1688980957
transform 1 0 35604 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2278_
timestamp 1688980957
transform -1 0 36984 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2279_
timestamp 1688980957
transform 1 0 36708 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _2280_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2281_
timestamp 1688980957
transform -1 0 12972 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2282_
timestamp 1688980957
transform -1 0 8832 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2283_
timestamp 1688980957
transform -1 0 13064 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2284_
timestamp 1688980957
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2285_
timestamp 1688980957
transform -1 0 13340 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2286_
timestamp 1688980957
transform 1 0 12972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2287_
timestamp 1688980957
transform -1 0 13156 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2288_
timestamp 1688980957
transform 1 0 1748 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2289_
timestamp 1688980957
transform 1 0 36616 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2290_
timestamp 1688980957
transform -1 0 37628 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _2291_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2292_
timestamp 1688980957
transform 1 0 1656 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2293_
timestamp 1688980957
transform 1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2294_
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2295_
timestamp 1688980957
transform -1 0 12972 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2296_
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2297_
timestamp 1688980957
transform 1 0 5796 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2298_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2299_
timestamp 1688980957
transform -1 0 5060 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2300_
timestamp 1688980957
transform 1 0 3864 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2301_
timestamp 1688980957
transform 1 0 7176 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2302_
timestamp 1688980957
transform -1 0 17572 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2303_
timestamp 1688980957
transform 1 0 2760 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2304_
timestamp 1688980957
transform 1 0 2944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2305_
timestamp 1688980957
transform 1 0 3864 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2306_
timestamp 1688980957
transform -1 0 9660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2307_
timestamp 1688980957
transform 1 0 3036 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2308_
timestamp 1688980957
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2309_
timestamp 1688980957
transform 1 0 5704 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2310_
timestamp 1688980957
transform -1 0 23000 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2311_
timestamp 1688980957
transform 1 0 17388 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2312_
timestamp 1688980957
transform -1 0 17664 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2313_
timestamp 1688980957
transform -1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2314_
timestamp 1688980957
transform 1 0 2668 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2315_
timestamp 1688980957
transform 1 0 1564 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2316_
timestamp 1688980957
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2317_
timestamp 1688980957
transform 1 0 2760 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2318_
timestamp 1688980957
transform 1 0 2208 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2319_
timestamp 1688980957
transform 1 0 5244 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2320_
timestamp 1688980957
transform -1 0 22908 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2321_
timestamp 1688980957
transform 1 0 7820 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2322_
timestamp 1688980957
transform -1 0 25392 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2323_
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2324_
timestamp 1688980957
transform -1 0 13064 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2325_
timestamp 1688980957
transform 1 0 4968 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2326_
timestamp 1688980957
transform 1 0 5428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2327_
timestamp 1688980957
transform -1 0 6348 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2328_
timestamp 1688980957
transform 1 0 2116 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2329_
timestamp 1688980957
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2330_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27416 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2331_
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2332_
timestamp 1688980957
transform -1 0 25300 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2333_
timestamp 1688980957
transform 1 0 18308 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2334_
timestamp 1688980957
transform -1 0 25392 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2335_
timestamp 1688980957
transform 1 0 1748 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2336_
timestamp 1688980957
transform 1 0 27232 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2337_
timestamp 1688980957
transform -1 0 37444 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2338_
timestamp 1688980957
transform -1 0 25852 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2339_
timestamp 1688980957
transform 1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2340_
timestamp 1688980957
transform 1 0 27508 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2341_
timestamp 1688980957
transform -1 0 34960 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2342_
timestamp 1688980957
transform 1 0 27968 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2343_
timestamp 1688980957
transform -1 0 32292 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2344_
timestamp 1688980957
transform -1 0 26220 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2345_
timestamp 1688980957
transform 1 0 4968 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2346_
timestamp 1688980957
transform -1 0 25760 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2347_
timestamp 1688980957
transform 1 0 12328 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2348_
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2349_
timestamp 1688980957
transform -1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2350_
timestamp 1688980957
transform 1 0 8188 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2351_
timestamp 1688980957
transform 1 0 9108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2352_
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2353_
timestamp 1688980957
transform 1 0 6440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2354_
timestamp 1688980957
transform 1 0 7084 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2355_
timestamp 1688980957
transform 1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2356_
timestamp 1688980957
transform 1 0 6624 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2357_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2358_
timestamp 1688980957
transform 1 0 6440 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2359_
timestamp 1688980957
transform 1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2360_
timestamp 1688980957
transform 1 0 9384 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2361_
timestamp 1688980957
transform 1 0 7176 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2362_
timestamp 1688980957
transform 1 0 6900 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2363_
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2364_
timestamp 1688980957
transform 1 0 8004 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2365_
timestamp 1688980957
transform 1 0 6900 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2366_
timestamp 1688980957
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2367_
timestamp 1688980957
transform 1 0 6532 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2368_
timestamp 1688980957
transform -1 0 6256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2369_
timestamp 1688980957
transform 1 0 7176 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2370_
timestamp 1688980957
transform 1 0 6992 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2371_
timestamp 1688980957
transform -1 0 13984 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2372_
timestamp 1688980957
transform -1 0 13156 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2373_
timestamp 1688980957
transform 1 0 11500 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2374_
timestamp 1688980957
transform -1 0 10948 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2375_
timestamp 1688980957
transform -1 0 13524 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2376_
timestamp 1688980957
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2377_
timestamp 1688980957
transform 1 0 15088 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2378_
timestamp 1688980957
transform -1 0 14996 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2379_
timestamp 1688980957
transform 1 0 12420 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2380_
timestamp 1688980957
transform -1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2381_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2382_
timestamp 1688980957
transform 1 0 10304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2383_
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2384_
timestamp 1688980957
transform -1 0 13984 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2385_
timestamp 1688980957
transform 1 0 11776 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2386_
timestamp 1688980957
transform -1 0 11684 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2387_
timestamp 1688980957
transform -1 0 13616 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2388_
timestamp 1688980957
transform 1 0 13616 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2389_
timestamp 1688980957
transform 1 0 9108 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2390_
timestamp 1688980957
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2391_
timestamp 1688980957
transform 1 0 15364 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2392_
timestamp 1688980957
transform -1 0 15732 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2393_
timestamp 1688980957
transform -1 0 16008 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2394_
timestamp 1688980957
transform 1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2395_
timestamp 1688980957
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2396_
timestamp 1688980957
transform -1 0 13432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2397_
timestamp 1688980957
transform 1 0 10304 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2398_
timestamp 1688980957
transform -1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2399_
timestamp 1688980957
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2400_
timestamp 1688980957
transform -1 0 15824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2401_
timestamp 1688980957
transform 1 0 10304 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2402_
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2403_
timestamp 1688980957
transform 1 0 9752 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2404_
timestamp 1688980957
transform 1 0 9476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2405_
timestamp 1688980957
transform 1 0 16192 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2406_
timestamp 1688980957
transform -1 0 30452 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2407__8
timestamp 1688980957
transform 1 0 10488 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2408__9
timestamp 1688980957
transform -1 0 7360 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2409__10
timestamp 1688980957
transform -1 0 6992 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2410__11
timestamp 1688980957
transform -1 0 4600 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2411__12
timestamp 1688980957
transform -1 0 6164 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2412__13
timestamp 1688980957
transform 1 0 3956 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2413__14
timestamp 1688980957
transform -1 0 9200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2414__15
timestamp 1688980957
transform 1 0 4508 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2415__16
timestamp 1688980957
transform -1 0 7636 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2416__17
timestamp 1688980957
transform 1 0 6624 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2417__18
timestamp 1688980957
transform -1 0 8372 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2418__19
timestamp 1688980957
transform -1 0 8188 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2419__20
timestamp 1688980957
transform -1 0 4232 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2420__21
timestamp 1688980957
transform 1 0 4048 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2421__22
timestamp 1688980957
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2422__23
timestamp 1688980957
transform 1 0 20148 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2423__24
timestamp 1688980957
transform -1 0 25944 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2424__25
timestamp 1688980957
transform 1 0 30360 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2425__26
timestamp 1688980957
transform 1 0 30728 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2426_
timestamp 1688980957
transform -1 0 34040 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2427__27
timestamp 1688980957
transform 1 0 34960 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2428__28
timestamp 1688980957
transform -1 0 35052 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2429__29
timestamp 1688980957
transform -1 0 31556 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2430__30
timestamp 1688980957
transform -1 0 27784 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2431__31
timestamp 1688980957
transform -1 0 32660 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2432__32
timestamp 1688980957
transform -1 0 9200 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2433__33
timestamp 1688980957
transform 1 0 5704 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2434__34
timestamp 1688980957
transform 1 0 9476 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2435__35
timestamp 1688980957
transform 1 0 5612 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2436__36
timestamp 1688980957
transform -1 0 4416 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2437__37
timestamp 1688980957
transform 1 0 4692 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2438__38
timestamp 1688980957
transform -1 0 13432 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2439__39
timestamp 1688980957
transform 1 0 21528 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2440__40
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2441__41
timestamp 1688980957
transform -1 0 33028 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2442__42
timestamp 1688980957
transform -1 0 33764 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2443__43
timestamp 1688980957
transform -1 0 34960 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2444__44
timestamp 1688980957
transform -1 0 32016 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2445__45
timestamp 1688980957
transform -1 0 27968 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2446_
timestamp 1688980957
transform -1 0 27048 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2447__46
timestamp 1688980957
transform 1 0 25024 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2448__47
timestamp 1688980957
transform 1 0 29624 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2449__48
timestamp 1688980957
transform -1 0 10488 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2450__49
timestamp 1688980957
transform -1 0 9568 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2451__50
timestamp 1688980957
transform 1 0 9936 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2452__51
timestamp 1688980957
transform 1 0 9200 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2453__52
timestamp 1688980957
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2454__53
timestamp 1688980957
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2455__54
timestamp 1688980957
transform 1 0 9016 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2456__55
timestamp 1688980957
transform 1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2457__56
timestamp 1688980957
transform -1 0 27968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2458__57
timestamp 1688980957
transform -1 0 28980 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2459__58
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2460__59
timestamp 1688980957
transform -1 0 27508 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2461__60
timestamp 1688980957
transform -1 0 29440 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2462__61
timestamp 1688980957
transform -1 0 28060 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2463__62
timestamp 1688980957
transform -1 0 27784 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2464__63
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2465__64
timestamp 1688980957
transform -1 0 29256 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2466__1
timestamp 1688980957
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2467__2
timestamp 1688980957
transform 1 0 35144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2468__3
timestamp 1688980957
transform -1 0 35144 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2469__4
timestamp 1688980957
transform -1 0 35144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2470__5
timestamp 1688980957
transform -1 0 30544 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2471__6
timestamp 1688980957
transform -1 0 27324 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2472__7
timestamp 1688980957
transform 1 0 34316 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2473_
timestamp 1688980957
transform 1 0 17480 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2474_
timestamp 1688980957
transform 1 0 18676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2475_
timestamp 1688980957
transform -1 0 10672 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2476_
timestamp 1688980957
transform -1 0 19136 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2477_
timestamp 1688980957
transform 1 0 10120 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2478_
timestamp 1688980957
transform -1 0 11408 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2479_
timestamp 1688980957
transform -1 0 12972 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2480_
timestamp 1688980957
transform -1 0 12512 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2481_
timestamp 1688980957
transform -1 0 13248 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2482_
timestamp 1688980957
transform -1 0 11316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2483_
timestamp 1688980957
transform -1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2484_
timestamp 1688980957
transform 1 0 11316 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2485_
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2486_
timestamp 1688980957
transform -1 0 12604 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2487_
timestamp 1688980957
transform -1 0 13064 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _2488_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12328 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _2489_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2490_
timestamp 1688980957
transform 1 0 11500 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _2491_
timestamp 1688980957
transform -1 0 12052 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2492_
timestamp 1688980957
transform 1 0 10304 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _2493_
timestamp 1688980957
transform 1 0 16008 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _2494_
timestamp 1688980957
transform -1 0 12696 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2495_
timestamp 1688980957
transform -1 0 11040 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2496_
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  _2497_
timestamp 1688980957
transform 1 0 13340 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _2498_
timestamp 1688980957
transform 1 0 8004 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2499_
timestamp 1688980957
transform 1 0 7636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2500_
timestamp 1688980957
transform 1 0 17572 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2501_
timestamp 1688980957
transform -1 0 17572 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2502_
timestamp 1688980957
transform -1 0 6992 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2503_
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2504_
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2505_
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2506_
timestamp 1688980957
transform 1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2507_
timestamp 1688980957
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2508_
timestamp 1688980957
transform -1 0 6808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2509_
timestamp 1688980957
transform 1 0 5612 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2510_
timestamp 1688980957
transform 1 0 5060 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2511_
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2512_
timestamp 1688980957
transform 1 0 3220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2513_
timestamp 1688980957
transform 1 0 13064 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2514_
timestamp 1688980957
transform -1 0 6164 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2515_
timestamp 1688980957
transform -1 0 6256 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2516_
timestamp 1688980957
transform -1 0 6256 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2517_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2518_
timestamp 1688980957
transform 1 0 5152 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2519_
timestamp 1688980957
transform 1 0 4600 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2520_
timestamp 1688980957
transform 1 0 10580 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2521_
timestamp 1688980957
transform 1 0 3128 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2522_
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2523_
timestamp 1688980957
transform 1 0 2300 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2524_
timestamp 1688980957
transform 1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2525_
timestamp 1688980957
transform 1 0 22172 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2526_
timestamp 1688980957
transform 1 0 17572 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2527_
timestamp 1688980957
transform -1 0 4232 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2528_
timestamp 1688980957
transform 1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2529_
timestamp 1688980957
transform 1 0 4416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2530_
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2531_
timestamp 1688980957
transform 1 0 2576 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2532_
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2533_
timestamp 1688980957
transform 1 0 10948 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2534_
timestamp 1688980957
transform 1 0 4508 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2535_
timestamp 1688980957
transform -1 0 3680 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2536_
timestamp 1688980957
transform 1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2537_
timestamp 1688980957
transform 1 0 3680 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2538_
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2539_
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2540_
timestamp 1688980957
transform 1 0 11868 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2541_
timestamp 1688980957
transform 1 0 4416 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2542_
timestamp 1688980957
transform 1 0 5152 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2543_
timestamp 1688980957
transform 1 0 4508 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2544_
timestamp 1688980957
transform 1 0 4232 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2545_
timestamp 1688980957
transform -1 0 4324 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2546_
timestamp 1688980957
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2547_
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _2548_
timestamp 1688980957
transform -1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2549_
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2550_
timestamp 1688980957
transform 1 0 2300 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2551_
timestamp 1688980957
transform 1 0 2024 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2552_
timestamp 1688980957
transform 1 0 3312 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2553_
timestamp 1688980957
transform 1 0 3772 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2554_
timestamp 1688980957
transform 1 0 3496 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2555_
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2556_
timestamp 1688980957
transform 1 0 2392 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2557_
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2558_
timestamp 1688980957
transform 1 0 3864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2559_
timestamp 1688980957
transform -1 0 3864 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2560_
timestamp 1688980957
transform 1 0 2944 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2561_
timestamp 1688980957
transform 1 0 2300 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2562_
timestamp 1688980957
transform 1 0 1748 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2563_
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2564_
timestamp 1688980957
transform 1 0 4232 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2565_
timestamp 1688980957
transform -1 0 4416 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2566_
timestamp 1688980957
transform 1 0 4048 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2567_
timestamp 1688980957
transform 1 0 3220 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2568_
timestamp 1688980957
transform 1 0 1748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2569_
timestamp 1688980957
transform 1 0 6716 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2570_
timestamp 1688980957
transform 1 0 7728 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2571_
timestamp 1688980957
transform 1 0 6992 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2572_
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2573_
timestamp 1688980957
transform 1 0 5704 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2574_
timestamp 1688980957
transform -1 0 6716 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2575_
timestamp 1688980957
transform -1 0 5704 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2576_
timestamp 1688980957
transform 1 0 5704 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2577_
timestamp 1688980957
transform 1 0 4968 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2578_
timestamp 1688980957
transform 1 0 4324 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2579_
timestamp 1688980957
transform 1 0 3864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2580_
timestamp 1688980957
transform -1 0 5796 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2581_
timestamp 1688980957
transform -1 0 5520 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2582_
timestamp 1688980957
transform 1 0 4232 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2583_
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2584_
timestamp 1688980957
transform 1 0 2852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2585_
timestamp 1688980957
transform 1 0 4508 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2586_
timestamp 1688980957
transform -1 0 6624 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2587_
timestamp 1688980957
transform 1 0 5152 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2588_
timestamp 1688980957
transform 1 0 4692 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2589_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2590_
timestamp 1688980957
transform 1 0 6900 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2591_
timestamp 1688980957
transform 1 0 8004 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2592_
timestamp 1688980957
transform 1 0 5060 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2593_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6164 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2594_
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2595_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2596_
timestamp 1688980957
transform 1 0 6532 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2597_
timestamp 1688980957
transform 1 0 7544 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2598_
timestamp 1688980957
transform 1 0 6072 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2599_
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2600_
timestamp 1688980957
transform 1 0 6624 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2601_
timestamp 1688980957
transform 1 0 10948 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2602_
timestamp 1688980957
transform 1 0 11868 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2603_
timestamp 1688980957
transform 1 0 15088 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2604_
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2605_
timestamp 1688980957
transform 1 0 9844 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2606_
timestamp 1688980957
transform 1 0 13892 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2607_
timestamp 1688980957
transform 1 0 11684 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2608_
timestamp 1688980957
transform 1 0 13156 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2609_
timestamp 1688980957
transform 1 0 8280 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2610_
timestamp 1688980957
transform 1 0 15456 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2611_
timestamp 1688980957
transform 1 0 15732 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2612_
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2613_
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2614_
timestamp 1688980957
transform 1 0 15824 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2615_
timestamp 1688980957
transform 1 0 9752 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2616_
timestamp 1688980957
transform 1 0 9108 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2617_
timestamp 1688980957
transform 1 0 10764 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2618_
timestamp 1688980957
transform 1 0 6992 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2619_
timestamp 1688980957
transform 1 0 6624 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2620_
timestamp 1688980957
transform 1 0 4232 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2621_
timestamp 1688980957
transform 1 0 6164 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2622_
timestamp 1688980957
transform 1 0 4232 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2623_
timestamp 1688980957
transform 1 0 8648 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2624_
timestamp 1688980957
transform 1 0 4784 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2625_
timestamp 1688980957
transform 1 0 7268 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2626_
timestamp 1688980957
transform 1 0 6900 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2627_
timestamp 1688980957
transform 1 0 7636 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2628_
timestamp 1688980957
transform 1 0 7820 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2629_
timestamp 1688980957
transform 1 0 3864 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2630_
timestamp 1688980957
transform 1 0 4324 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2631_
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2632_
timestamp 1688980957
transform 1 0 20424 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2633_
timestamp 1688980957
transform 1 0 25576 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2634_
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2635_
timestamp 1688980957
transform 1 0 31004 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2636_
timestamp 1688980957
transform 1 0 34500 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2637_
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2638_
timestamp 1688980957
transform 1 0 31188 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2639_
timestamp 1688980957
transform 1 0 27416 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2640_
timestamp 1688980957
transform 1 0 32292 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2641_
timestamp 1688980957
transform 1 0 8648 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2642_
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2643_
timestamp 1688980957
transform 1 0 9752 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2644_
timestamp 1688980957
transform 1 0 5888 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2645_
timestamp 1688980957
transform 1 0 4048 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2646_
timestamp 1688980957
transform 1 0 4968 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2647_
timestamp 1688980957
transform -1 0 13156 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2648_
timestamp 1688980957
transform 1 0 21804 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2649_
timestamp 1688980957
transform 1 0 25760 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2650_
timestamp 1688980957
transform 1 0 32660 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2651_
timestamp 1688980957
transform 1 0 33396 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2652_
timestamp 1688980957
transform -1 0 34500 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2653_
timestamp 1688980957
transform 1 0 31740 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2654_
timestamp 1688980957
transform 1 0 27508 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2655_
timestamp 1688980957
transform 1 0 25300 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2656_
timestamp 1688980957
transform 1 0 29900 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2657_
timestamp 1688980957
transform 1 0 10120 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2658_
timestamp 1688980957
transform 1 0 9200 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2659_
timestamp 1688980957
transform 1 0 10212 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2660_
timestamp 1688980957
transform 1 0 9476 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2661_
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2662_
timestamp 1688980957
transform 1 0 8924 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2663_
timestamp 1688980957
transform 1 0 9292 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2664_
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2665_
timestamp 1688980957
transform 1 0 27508 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2666_
timestamp 1688980957
transform 1 0 28612 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2667_
timestamp 1688980957
transform 1 0 29440 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2668_
timestamp 1688980957
transform 1 0 27232 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2669_
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2670_
timestamp 1688980957
transform 1 0 27692 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2671_
timestamp 1688980957
transform 1 0 27232 0 1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2672_
timestamp 1688980957
transform 1 0 29072 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2673_
timestamp 1688980957
transform 1 0 28888 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2674_
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2675_
timestamp 1688980957
transform 1 0 34960 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2676_
timestamp 1688980957
transform 1 0 34776 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2677_
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2678_
timestamp 1688980957
transform 1 0 29900 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2679_
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2680_
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2681_
timestamp 1688980957
transform 1 0 6900 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2682_
timestamp 1688980957
transform 1 0 4232 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2683_
timestamp 1688980957
transform 1 0 2576 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2684_
timestamp 1688980957
transform 1 0 4048 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2685_
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2686_
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2687_
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2688_
timestamp 1688980957
transform 1 0 3956 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2689_
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2690_
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2691_
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2692_
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2693_
timestamp 1688980957
transform 1 0 5244 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2694_
timestamp 1688980957
transform 1 0 3312 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2695_
timestamp 1688980957
transform 1 0 1840 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2696_
timestamp 1688980957
transform 1 0 4140 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2697_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17572 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2698_
timestamp 1688980957
transform 1 0 13432 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2699_
timestamp 1688980957
transform 1 0 10672 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2700_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2701_
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2702_
timestamp 1688980957
transform 1 0 9384 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0514_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30912 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0515_
timestamp 1688980957
transform -1 0 19136 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0516_
timestamp 1688980957
transform -1 0 21344 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0517_
timestamp 1688980957
transform -1 0 21344 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0514_
timestamp 1688980957
transform 1 0 31188 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0515_
timestamp 1688980957
transform -1 0 11408 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0516_
timestamp 1688980957
transform -1 0 14812 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0517_
timestamp 1688980957
transform -1 0 14812 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0514_
timestamp 1688980957
transform -1 0 30452 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0515_
timestamp 1688980957
transform 1 0 20792 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0516_
timestamp 1688980957
transform 1 0 23368 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0517_
timestamp 1688980957
transform 1 0 23368 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1688980957
transform 1 0 7820 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1688980957
transform -1 0 4416 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1688980957
transform 1 0 9476 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  fanout57
timestamp 1688980957
transform 1 0 7820 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout58
timestamp 1688980957
transform -1 0 3404 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout59
timestamp 1688980957
transform -1 0 9200 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout60
timestamp 1688980957
transform 1 0 7176 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout61
timestamp 1688980957
transform -1 0 8832 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  fanout62
timestamp 1688980957
transform 1 0 28336 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout63
timestamp 1688980957
transform 1 0 20240 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_97 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_105
timestamp 1688980957
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_125 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_135
timestamp 1688980957
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_149
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_156
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_184
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_205
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_217
timestamp 1688980957
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_287
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_299
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_399
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_10
timestamp 1688980957
transform 1 0 2024 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_121
timestamp 1688980957
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_132
timestamp 1688980957
transform 1 0 13248 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_153
timestamp 1688980957
transform 1 0 15180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_165
timestamp 1688980957
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_178
timestamp 1688980957
transform 1 0 17480 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_190
timestamp 1688980957
transform 1 0 18584 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_202
timestamp 1688980957
transform 1 0 19688 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_206
timestamp 1688980957
transform 1 0 20056 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_218
timestamp 1688980957
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_95
timestamp 1688980957
transform 1 0 9844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_107
timestamp 1688980957
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_143
timestamp 1688980957
transform 1 0 14260 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_147
timestamp 1688980957
transform 1 0 14628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_159
timestamp 1688980957
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_257
timestamp 1688980957
transform 1 0 24748 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_265
timestamp 1688980957
transform 1 0 25484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_277
timestamp 1688980957
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_289
timestamp 1688980957
transform 1 0 27692 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_9
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_21
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_93
timestamp 1688980957
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_100
timestamp 1688980957
transform 1 0 10304 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_125
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_137
timestamp 1688980957
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_169
timestamp 1688980957
transform 1 0 16652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_181
timestamp 1688980957
transform 1 0 17756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_204
timestamp 1688980957
transform 1 0 19872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_210
timestamp 1688980957
transform 1 0 20424 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_244
timestamp 1688980957
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_318
timestamp 1688980957
transform 1 0 30360 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_330
timestamp 1688980957
transform 1 0 31464 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_342
timestamp 1688980957
transform 1 0 32568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_354
timestamp 1688980957
transform 1 0 33672 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_362
timestamp 1688980957
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_61
timestamp 1688980957
transform 1 0 6716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_73
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_85
timestamp 1688980957
transform 1 0 8924 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_101
timestamp 1688980957
transform 1 0 10396 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_110
timestamp 1688980957
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_154
timestamp 1688980957
transform 1 0 15272 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_158
timestamp 1688980957
transform 1 0 15640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_177
timestamp 1688980957
transform 1 0 17388 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_189
timestamp 1688980957
transform 1 0 18492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_197
timestamp 1688980957
transform 1 0 19228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_206
timestamp 1688980957
transform 1 0 20056 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_214
timestamp 1688980957
transform 1 0 20792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_220
timestamp 1688980957
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_241
timestamp 1688980957
transform 1 0 23276 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_246
timestamp 1688980957
transform 1 0 23736 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_258
timestamp 1688980957
transform 1 0 24840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_270
timestamp 1688980957
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 1688980957
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_292
timestamp 1688980957
transform 1 0 27968 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_331
timestamp 1688980957
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_106
timestamp 1688980957
transform 1 0 10856 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_129
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_179
timestamp 1688980957
transform 1 0 17572 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_191
timestamp 1688980957
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_205
timestamp 1688980957
transform 1 0 19964 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_213
timestamp 1688980957
transform 1 0 20700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_225
timestamp 1688980957
transform 1 0 21804 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_248
timestamp 1688980957
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_261
timestamp 1688980957
transform 1 0 25116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_273
timestamp 1688980957
transform 1 0 26220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_285
timestamp 1688980957
transform 1 0 27324 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_297
timestamp 1688980957
transform 1 0 28428 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_305
timestamp 1688980957
transform 1 0 29164 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_320
timestamp 1688980957
transform 1 0 30544 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_340
timestamp 1688980957
transform 1 0 32384 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_352
timestamp 1688980957
transform 1 0 33488 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_42
timestamp 1688980957
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1688980957
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_94
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_130
timestamp 1688980957
transform 1 0 13064 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_160
timestamp 1688980957
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_198
timestamp 1688980957
transform 1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_239
timestamp 1688980957
transform 1 0 23092 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_247
timestamp 1688980957
transform 1 0 23828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_254
timestamp 1688980957
transform 1 0 24472 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_262
timestamp 1688980957
transform 1 0 25208 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_267
timestamp 1688980957
transform 1 0 25668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_296
timestamp 1688980957
transform 1 0 28336 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_308
timestamp 1688980957
transform 1 0 29440 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_320
timestamp 1688980957
transform 1 0 30544 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_332
timestamp 1688980957
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_345
timestamp 1688980957
transform 1 0 32844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_357
timestamp 1688980957
transform 1 0 33948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_369
timestamp 1688980957
transform 1 0 35052 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_381
timestamp 1688980957
transform 1 0 36156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_389
timestamp 1688980957
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_33
timestamp 1688980957
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_54
timestamp 1688980957
transform 1 0 6072 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_66
timestamp 1688980957
transform 1 0 7176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_78
timestamp 1688980957
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_88
timestamp 1688980957
transform 1 0 9200 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_100
timestamp 1688980957
transform 1 0 10304 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_112
timestamp 1688980957
transform 1 0 11408 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_120
timestamp 1688980957
transform 1 0 12144 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_129
timestamp 1688980957
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1688980957
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_145
timestamp 1688980957
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_154
timestamp 1688980957
transform 1 0 15272 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_176
timestamp 1688980957
transform 1 0 17296 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_203
timestamp 1688980957
transform 1 0 19780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_211
timestamp 1688980957
transform 1 0 20516 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_217
timestamp 1688980957
transform 1 0 21068 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_224
timestamp 1688980957
transform 1 0 21712 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_236
timestamp 1688980957
transform 1 0 22816 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_248
timestamp 1688980957
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_268
timestamp 1688980957
transform 1 0 25760 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_278
timestamp 1688980957
transform 1 0 26680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_285
timestamp 1688980957
transform 1 0 27324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_302
timestamp 1688980957
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_325
timestamp 1688980957
transform 1 0 31004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_329
timestamp 1688980957
transform 1 0 31372 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_338
timestamp 1688980957
transform 1 0 32200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_354
timestamp 1688980957
transform 1 0 33672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_362
timestamp 1688980957
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_7
timestamp 1688980957
transform 1 0 1748 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_36
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_64
timestamp 1688980957
transform 1 0 6992 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_70
timestamp 1688980957
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_74
timestamp 1688980957
transform 1 0 7912 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_86
timestamp 1688980957
transform 1 0 9016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1688980957
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_133
timestamp 1688980957
transform 1 0 13340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_152
timestamp 1688980957
transform 1 0 15088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_159
timestamp 1688980957
transform 1 0 15732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_184
timestamp 1688980957
transform 1 0 18032 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_192
timestamp 1688980957
transform 1 0 18768 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_199
timestamp 1688980957
transform 1 0 19412 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_210
timestamp 1688980957
transform 1 0 20424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_219
timestamp 1688980957
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_232
timestamp 1688980957
transform 1 0 22448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_241
timestamp 1688980957
transform 1 0 23276 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_267
timestamp 1688980957
transform 1 0 25668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_278
timestamp 1688980957
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_287
timestamp 1688980957
transform 1 0 27508 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_318
timestamp 1688980957
transform 1 0 30360 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_52
timestamp 1688980957
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_96
timestamp 1688980957
transform 1 0 9936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_100
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_164
timestamp 1688980957
transform 1 0 16192 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_172
timestamp 1688980957
transform 1 0 16928 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_182
timestamp 1688980957
transform 1 0 17848 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1688980957
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_201
timestamp 1688980957
transform 1 0 19596 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_205
timestamp 1688980957
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_313
timestamp 1688980957
transform 1 0 29900 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_323
timestamp 1688980957
transform 1 0 30820 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_335
timestamp 1688980957
transform 1 0 31924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_347
timestamp 1688980957
transform 1 0 33028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_359
timestamp 1688980957
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_26
timestamp 1688980957
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_38
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_42
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_62
timestamp 1688980957
transform 1 0 6808 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_70
timestamp 1688980957
transform 1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_154
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1688980957
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_180
timestamp 1688980957
transform 1 0 17664 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_195
timestamp 1688980957
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_199
timestamp 1688980957
transform 1 0 19412 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_204
timestamp 1688980957
transform 1 0 19872 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_216
timestamp 1688980957
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_231
timestamp 1688980957
transform 1 0 22356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_246
timestamp 1688980957
transform 1 0 23736 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_254
timestamp 1688980957
transform 1 0 24472 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_264
timestamp 1688980957
transform 1 0 25392 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_276
timestamp 1688980957
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_290
timestamp 1688980957
transform 1 0 27784 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_308
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_320
timestamp 1688980957
transform 1 0 30544 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_326
timestamp 1688980957
transform 1 0 31096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_343
timestamp 1688980957
transform 1 0 32660 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_351
timestamp 1688980957
transform 1 0 33396 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_363
timestamp 1688980957
transform 1 0 34500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_375
timestamp 1688980957
transform 1 0 35604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_387
timestamp 1688980957
transform 1 0 36708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 1688980957
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_43
timestamp 1688980957
transform 1 0 5060 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_56
timestamp 1688980957
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_68
timestamp 1688980957
transform 1 0 7360 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_74
timestamp 1688980957
transform 1 0 7912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_93
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_114
timestamp 1688980957
transform 1 0 11592 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1688980957
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_149
timestamp 1688980957
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_179
timestamp 1688980957
transform 1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_192
timestamp 1688980957
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_206
timestamp 1688980957
transform 1 0 20056 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_216
timestamp 1688980957
transform 1 0 20976 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_228
timestamp 1688980957
transform 1 0 22080 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1688980957
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_261
timestamp 1688980957
transform 1 0 25116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_293
timestamp 1688980957
transform 1 0 28060 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_319
timestamp 1688980957
transform 1 0 30452 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_325
timestamp 1688980957
transform 1 0 31004 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_339
timestamp 1688980957
transform 1 0 32292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_353
timestamp 1688980957
transform 1 0 33580 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_361
timestamp 1688980957
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_19
timestamp 1688980957
transform 1 0 2852 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_28
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_40
timestamp 1688980957
transform 1 0 4784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_52
timestamp 1688980957
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_65
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_79
timestamp 1688980957
transform 1 0 8372 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_83
timestamp 1688980957
transform 1 0 8740 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_95
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_129
timestamp 1688980957
transform 1 0 12972 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_139
timestamp 1688980957
transform 1 0 13892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_151
timestamp 1688980957
transform 1 0 14996 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 1688980957
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_178
timestamp 1688980957
transform 1 0 17480 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_200
timestamp 1688980957
transform 1 0 19504 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_208
timestamp 1688980957
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_220
timestamp 1688980957
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_231
timestamp 1688980957
transform 1 0 22356 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_240
timestamp 1688980957
transform 1 0 23184 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_248
timestamp 1688980957
transform 1 0 23920 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_260
timestamp 1688980957
transform 1 0 25024 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_268
timestamp 1688980957
transform 1 0 25760 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_289
timestamp 1688980957
transform 1 0 27692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_306
timestamp 1688980957
transform 1 0 29256 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_316
timestamp 1688980957
transform 1 0 30176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_344
timestamp 1688980957
transform 1 0 32752 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_350
timestamp 1688980957
transform 1 0 33304 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_362
timestamp 1688980957
transform 1 0 34408 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_374
timestamp 1688980957
transform 1 0 35512 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_386
timestamp 1688980957
transform 1 0 36616 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_23
timestamp 1688980957
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_37
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_56
timestamp 1688980957
transform 1 0 6256 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_68
timestamp 1688980957
transform 1 0 7360 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1688980957
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_92
timestamp 1688980957
transform 1 0 9568 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_104
timestamp 1688980957
transform 1 0 10672 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1688980957
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_192
timestamp 1688980957
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_203
timestamp 1688980957
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_207
timestamp 1688980957
transform 1 0 20148 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_227
timestamp 1688980957
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_235
timestamp 1688980957
transform 1 0 22724 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_247
timestamp 1688980957
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_289
timestamp 1688980957
transform 1 0 27692 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_305
timestamp 1688980957
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_324
timestamp 1688980957
transform 1 0 30912 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_336
timestamp 1688980957
transform 1 0 32016 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_345
timestamp 1688980957
transform 1 0 32844 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_351
timestamp 1688980957
transform 1 0 33396 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_360
timestamp 1688980957
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1688980957
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1688980957
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_10
timestamp 1688980957
transform 1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_29
timestamp 1688980957
transform 1 0 3772 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_52
timestamp 1688980957
transform 1 0 5888 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_71
timestamp 1688980957
transform 1 0 7636 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_79
timestamp 1688980957
transform 1 0 8372 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_101
timestamp 1688980957
transform 1 0 10396 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_162
timestamp 1688980957
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_179
timestamp 1688980957
transform 1 0 17572 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_202
timestamp 1688980957
transform 1 0 19688 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_209
timestamp 1688980957
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_213
timestamp 1688980957
transform 1 0 20700 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_233
timestamp 1688980957
transform 1 0 22540 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_243
timestamp 1688980957
transform 1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_256
timestamp 1688980957
transform 1 0 24656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_268
timestamp 1688980957
transform 1 0 25760 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_289
timestamp 1688980957
transform 1 0 27692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_304
timestamp 1688980957
transform 1 0 29072 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_316
timestamp 1688980957
transform 1 0 30176 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_320
timestamp 1688980957
transform 1 0 30544 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_332
timestamp 1688980957
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_347
timestamp 1688980957
transform 1 0 33028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_351
timestamp 1688980957
transform 1 0 33396 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_370
timestamp 1688980957
transform 1 0 35144 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_382
timestamp 1688980957
transform 1 0 36248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_390
timestamp 1688980957
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_23
timestamp 1688980957
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_38
timestamp 1688980957
transform 1 0 4600 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_55
timestamp 1688980957
transform 1 0 6164 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_67
timestamp 1688980957
transform 1 0 7268 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_92
timestamp 1688980957
transform 1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_117
timestamp 1688980957
transform 1 0 11868 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_132
timestamp 1688980957
transform 1 0 13248 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_136
timestamp 1688980957
transform 1 0 13616 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_150
timestamp 1688980957
transform 1 0 14904 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_156
timestamp 1688980957
transform 1 0 15456 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_180
timestamp 1688980957
transform 1 0 17664 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_193
timestamp 1688980957
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_217
timestamp 1688980957
transform 1 0 21068 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_241
timestamp 1688980957
transform 1 0 23276 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_247
timestamp 1688980957
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_261
timestamp 1688980957
transform 1 0 25116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_267
timestamp 1688980957
transform 1 0 25668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_298
timestamp 1688980957
transform 1 0 28520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_313
timestamp 1688980957
transform 1 0 29900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_350
timestamp 1688980957
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_362
timestamp 1688980957
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 1688980957
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_389
timestamp 1688980957
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_7
timestamp 1688980957
transform 1 0 1748 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_19
timestamp 1688980957
transform 1 0 2852 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_31
timestamp 1688980957
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_43
timestamp 1688980957
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_99
timestamp 1688980957
transform 1 0 10212 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1688980957
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_117
timestamp 1688980957
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_144
timestamp 1688980957
transform 1 0 14352 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_156
timestamp 1688980957
transform 1 0 15456 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1688980957
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_189
timestamp 1688980957
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_248
timestamp 1688980957
transform 1 0 23920 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_292
timestamp 1688980957
transform 1 0 27968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_304
timestamp 1688980957
transform 1 0 29072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_314
timestamp 1688980957
transform 1 0 29992 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_324
timestamp 1688980957
transform 1 0 30912 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_345
timestamp 1688980957
transform 1 0 32844 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_357
timestamp 1688980957
transform 1 0 33948 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_369
timestamp 1688980957
transform 1 0 35052 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_381
timestamp 1688980957
transform 1 0 36156 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_389
timestamp 1688980957
transform 1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_12
timestamp 1688980957
transform 1 0 2208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_25
timestamp 1688980957
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_38
timestamp 1688980957
transform 1 0 4600 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_50
timestamp 1688980957
transform 1 0 5704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_67
timestamp 1688980957
transform 1 0 7268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_93
timestamp 1688980957
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_99
timestamp 1688980957
transform 1 0 10212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_111
timestamp 1688980957
transform 1 0 11316 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_122
timestamp 1688980957
transform 1 0 12328 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_134
timestamp 1688980957
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_147
timestamp 1688980957
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_151
timestamp 1688980957
transform 1 0 14996 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_172
timestamp 1688980957
transform 1 0 16928 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_178
timestamp 1688980957
transform 1 0 17480 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_202
timestamp 1688980957
transform 1 0 19688 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_214
timestamp 1688980957
transform 1 0 20792 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_227
timestamp 1688980957
transform 1 0 21988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_235
timestamp 1688980957
transform 1 0 22724 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_247
timestamp 1688980957
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_261
timestamp 1688980957
transform 1 0 25116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_271
timestamp 1688980957
transform 1 0 26036 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_281
timestamp 1688980957
transform 1 0 26956 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_293
timestamp 1688980957
transform 1 0 28060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_305
timestamp 1688980957
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_345
timestamp 1688980957
transform 1 0 32844 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_356
timestamp 1688980957
transform 1 0 33856 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1688980957
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1688980957
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_23
timestamp 1688980957
transform 1 0 3220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_45
timestamp 1688980957
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_104
timestamp 1688980957
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_119
timestamp 1688980957
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_182
timestamp 1688980957
transform 1 0 17848 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_194
timestamp 1688980957
transform 1 0 18952 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_212
timestamp 1688980957
transform 1 0 20608 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_216
timestamp 1688980957
transform 1 0 20976 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_234
timestamp 1688980957
transform 1 0 22632 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_246
timestamp 1688980957
transform 1 0 23736 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_263
timestamp 1688980957
transform 1 0 25300 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_271
timestamp 1688980957
transform 1 0 26036 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_301
timestamp 1688980957
transform 1 0 28796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_308
timestamp 1688980957
transform 1 0 29440 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_316
timestamp 1688980957
transform 1 0 30176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_326
timestamp 1688980957
transform 1 0 31096 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1688980957
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_342
timestamp 1688980957
transform 1 0 32568 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1688980957
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 1688980957
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 1688980957
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1688980957
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_58
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_68
timestamp 1688980957
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_80
timestamp 1688980957
transform 1 0 8464 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_149
timestamp 1688980957
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_156
timestamp 1688980957
transform 1 0 15456 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_164
timestamp 1688980957
transform 1 0 16192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_172
timestamp 1688980957
transform 1 0 16928 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_180
timestamp 1688980957
transform 1 0 17664 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_184
timestamp 1688980957
transform 1 0 18032 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_201
timestamp 1688980957
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_215
timestamp 1688980957
transform 1 0 20884 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_225
timestamp 1688980957
transform 1 0 21804 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_246
timestamp 1688980957
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_258
timestamp 1688980957
transform 1 0 24840 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_266
timestamp 1688980957
transform 1 0 25576 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_287
timestamp 1688980957
transform 1 0 27508 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_301
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_312
timestamp 1688980957
transform 1 0 29808 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_324
timestamp 1688980957
transform 1 0 30912 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_336
timestamp 1688980957
transform 1 0 32016 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_340
timestamp 1688980957
transform 1 0 32384 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_359
timestamp 1688980957
transform 1 0 34132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1688980957
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 1688980957
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1688980957
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_12
timestamp 1688980957
transform 1 0 2208 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_24
timestamp 1688980957
transform 1 0 3312 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_36
timestamp 1688980957
transform 1 0 4416 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_48
timestamp 1688980957
transform 1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_77
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_83
timestamp 1688980957
transform 1 0 8740 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_95
timestamp 1688980957
transform 1 0 9844 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1688980957
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_143
timestamp 1688980957
transform 1 0 14260 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_176
timestamp 1688980957
transform 1 0 17296 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_186
timestamp 1688980957
transform 1 0 18216 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_198
timestamp 1688980957
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_285
timestamp 1688980957
transform 1 0 27324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_307
timestamp 1688980957
transform 1 0 29348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_315
timestamp 1688980957
transform 1 0 30084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_325
timestamp 1688980957
transform 1 0 31004 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_343
timestamp 1688980957
transform 1 0 32660 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_350
timestamp 1688980957
transform 1 0 33304 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_362
timestamp 1688980957
transform 1 0 34408 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_374
timestamp 1688980957
transform 1 0 35512 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_386
timestamp 1688980957
transform 1 0 36616 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_23
timestamp 1688980957
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_35
timestamp 1688980957
transform 1 0 4324 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_47
timestamp 1688980957
transform 1 0 5428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_70
timestamp 1688980957
transform 1 0 7544 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1688980957
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_93
timestamp 1688980957
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_118
timestamp 1688980957
transform 1 0 11960 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_135
timestamp 1688980957
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_160
timestamp 1688980957
transform 1 0 15824 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_171
timestamp 1688980957
transform 1 0 16836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_179
timestamp 1688980957
transform 1 0 17572 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_186
timestamp 1688980957
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_205
timestamp 1688980957
transform 1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_224
timestamp 1688980957
transform 1 0 21712 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_247
timestamp 1688980957
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1688980957
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_315
timestamp 1688980957
transform 1 0 30084 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_326
timestamp 1688980957
transform 1 0 31096 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_336
timestamp 1688980957
transform 1 0 32016 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_348
timestamp 1688980957
transform 1 0 33120 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_360
timestamp 1688980957
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1688980957
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1688980957
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_24
timestamp 1688980957
transform 1 0 3312 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_42
timestamp 1688980957
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1688980957
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_63
timestamp 1688980957
transform 1 0 6900 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_95
timestamp 1688980957
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_99
timestamp 1688980957
transform 1 0 10212 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_103
timestamp 1688980957
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_122
timestamp 1688980957
transform 1 0 12328 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_153
timestamp 1688980957
transform 1 0 15180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_160
timestamp 1688980957
transform 1 0 15824 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_187
timestamp 1688980957
transform 1 0 18308 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_203
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_212
timestamp 1688980957
transform 1 0 20608 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_230
timestamp 1688980957
transform 1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_242
timestamp 1688980957
transform 1 0 23368 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_254
timestamp 1688980957
transform 1 0 24472 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_262
timestamp 1688980957
transform 1 0 25208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_271
timestamp 1688980957
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_304
timestamp 1688980957
transform 1 0 29072 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_316
timestamp 1688980957
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_320
timestamp 1688980957
transform 1 0 30544 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_327
timestamp 1688980957
transform 1 0 31188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_352
timestamp 1688980957
transform 1 0 33488 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_362
timestamp 1688980957
transform 1 0 34408 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_374
timestamp 1688980957
transform 1 0 35512 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_386
timestamp 1688980957
transform 1 0 36616 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_9
timestamp 1688980957
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_21
timestamp 1688980957
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_43
timestamp 1688980957
transform 1 0 5060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_76
timestamp 1688980957
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_105
timestamp 1688980957
transform 1 0 10764 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_116
timestamp 1688980957
transform 1 0 11776 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_149
timestamp 1688980957
transform 1 0 14812 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_155
timestamp 1688980957
transform 1 0 15364 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_166
timestamp 1688980957
transform 1 0 16376 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_178
timestamp 1688980957
transform 1 0 17480 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_216
timestamp 1688980957
transform 1 0 20976 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_228
timestamp 1688980957
transform 1 0 22080 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_236
timestamp 1688980957
transform 1 0 22816 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_247
timestamp 1688980957
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_267
timestamp 1688980957
transform 1 0 25668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_279
timestamp 1688980957
transform 1 0 26772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_283
timestamp 1688980957
transform 1 0 27140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_291
timestamp 1688980957
transform 1 0 27876 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1688980957
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_322
timestamp 1688980957
transform 1 0 30728 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_335
timestamp 1688980957
transform 1 0 31924 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_352
timestamp 1688980957
transform 1 0 33488 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_379
timestamp 1688980957
transform 1 0 35972 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_391
timestamp 1688980957
transform 1 0 37076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_399
timestamp 1688980957
transform 1 0 37812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_23
timestamp 1688980957
transform 1 0 3220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_29
timestamp 1688980957
transform 1 0 3772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_35
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_43
timestamp 1688980957
transform 1 0 5060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1688980957
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_89
timestamp 1688980957
transform 1 0 9292 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_103
timestamp 1688980957
transform 1 0 10580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_126
timestamp 1688980957
transform 1 0 12696 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_138
timestamp 1688980957
transform 1 0 13800 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_176
timestamp 1688980957
transform 1 0 17296 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_197
timestamp 1688980957
transform 1 0 19228 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_205
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_214
timestamp 1688980957
transform 1 0 20792 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_222
timestamp 1688980957
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_233
timestamp 1688980957
transform 1 0 22540 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_243
timestamp 1688980957
transform 1 0 23460 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_249
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_277
timestamp 1688980957
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_288
timestamp 1688980957
transform 1 0 27600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_300
timestamp 1688980957
transform 1 0 28704 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_312
timestamp 1688980957
transform 1 0 29808 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_318
timestamp 1688980957
transform 1 0 30360 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_330
timestamp 1688980957
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_361
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_371
timestamp 1688980957
transform 1 0 35236 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_383
timestamp 1688980957
transform 1 0 36340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1688980957
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_393
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_22
timestamp 1688980957
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_40
timestamp 1688980957
transform 1 0 4784 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_52
timestamp 1688980957
transform 1 0 5888 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_64
timestamp 1688980957
transform 1 0 6992 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_76
timestamp 1688980957
transform 1 0 8096 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_107
timestamp 1688980957
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_119
timestamp 1688980957
transform 1 0 12052 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_131
timestamp 1688980957
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_176
timestamp 1688980957
transform 1 0 17296 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_205
timestamp 1688980957
transform 1 0 19964 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_238
timestamp 1688980957
transform 1 0 23000 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_249
timestamp 1688980957
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_261
timestamp 1688980957
transform 1 0 25116 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_267
timestamp 1688980957
transform 1 0 25668 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_276
timestamp 1688980957
transform 1 0 26496 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_288
timestamp 1688980957
transform 1 0 27600 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_300
timestamp 1688980957
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_313
timestamp 1688980957
transform 1 0 29900 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_317
timestamp 1688980957
transform 1 0 30268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_323
timestamp 1688980957
transform 1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_330
timestamp 1688980957
transform 1 0 31464 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_336
timestamp 1688980957
transform 1 0 32016 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_342
timestamp 1688980957
transform 1 0 32568 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_354
timestamp 1688980957
transform 1 0 33672 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_378
timestamp 1688980957
transform 1 0 35880 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_390
timestamp 1688980957
transform 1 0 36984 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_398
timestamp 1688980957
transform 1 0 37720 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_26
timestamp 1688980957
transform 1 0 3496 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_46
timestamp 1688980957
transform 1 0 5336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_62
timestamp 1688980957
transform 1 0 6808 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_72
timestamp 1688980957
transform 1 0 7728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_84
timestamp 1688980957
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_90
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_104
timestamp 1688980957
transform 1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_117
timestamp 1688980957
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_124
timestamp 1688980957
transform 1 0 12512 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_136
timestamp 1688980957
transform 1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_146
timestamp 1688980957
transform 1 0 14536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_158
timestamp 1688980957
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1688980957
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_174
timestamp 1688980957
transform 1 0 17112 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_186
timestamp 1688980957
transform 1 0 18216 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_198
timestamp 1688980957
transform 1 0 19320 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_245
timestamp 1688980957
transform 1 0 23644 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_257
timestamp 1688980957
transform 1 0 24748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_269
timestamp 1688980957
transform 1 0 25852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_277
timestamp 1688980957
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_289
timestamp 1688980957
transform 1 0 27692 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_301
timestamp 1688980957
transform 1 0 28796 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_310
timestamp 1688980957
transform 1 0 29624 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_322
timestamp 1688980957
transform 1 0 30728 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_330
timestamp 1688980957
transform 1 0 31464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_350
timestamp 1688980957
transform 1 0 33304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_354
timestamp 1688980957
transform 1 0 33672 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_360
timestamp 1688980957
transform 1 0 34224 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_371
timestamp 1688980957
transform 1 0 35236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_383
timestamp 1688980957
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_13
timestamp 1688980957
transform 1 0 2300 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_19
timestamp 1688980957
transform 1 0 2852 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_51
timestamp 1688980957
transform 1 0 5796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_78
timestamp 1688980957
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_94
timestamp 1688980957
transform 1 0 9752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_132
timestamp 1688980957
transform 1 0 13248 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_151
timestamp 1688980957
transform 1 0 14996 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_170
timestamp 1688980957
transform 1 0 16744 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_176
timestamp 1688980957
transform 1 0 17296 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_191
timestamp 1688980957
transform 1 0 18676 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_214
timestamp 1688980957
transform 1 0 20792 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_226
timestamp 1688980957
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_238
timestamp 1688980957
transform 1 0 23000 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_249
timestamp 1688980957
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_267
timestamp 1688980957
transform 1 0 25668 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_278
timestamp 1688980957
transform 1 0 26680 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_287
timestamp 1688980957
transform 1 0 27508 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_306
timestamp 1688980957
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_320
timestamp 1688980957
transform 1 0 30544 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_326
timestamp 1688980957
transform 1 0 31096 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_330
timestamp 1688980957
transform 1 0 31464 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_339
timestamp 1688980957
transform 1 0 32292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_351
timestamp 1688980957
transform 1 0 33396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_359
timestamp 1688980957
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 1688980957
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 1688980957
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_36
timestamp 1688980957
transform 1 0 4416 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_48
timestamp 1688980957
transform 1 0 5520 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_153
timestamp 1688980957
transform 1 0 15180 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_163
timestamp 1688980957
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_245
timestamp 1688980957
transform 1 0 23644 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_257
timestamp 1688980957
transform 1 0 24748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_274
timestamp 1688980957
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_289
timestamp 1688980957
transform 1 0 27692 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_295
timestamp 1688980957
transform 1 0 28244 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_307
timestamp 1688980957
transform 1 0 29348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_313
timestamp 1688980957
transform 1 0 29900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_324
timestamp 1688980957
transform 1 0 30912 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_373
timestamp 1688980957
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_385
timestamp 1688980957
transform 1 0 36524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_9
timestamp 1688980957
transform 1 0 1932 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1688980957
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_37
timestamp 1688980957
transform 1 0 4508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_42
timestamp 1688980957
transform 1 0 4968 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_48
timestamp 1688980957
transform 1 0 5520 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_57
timestamp 1688980957
transform 1 0 6348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_69
timestamp 1688980957
transform 1 0 7452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1688980957
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_147
timestamp 1688980957
transform 1 0 14628 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_159
timestamp 1688980957
transform 1 0 15732 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_171
timestamp 1688980957
transform 1 0 16836 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_191
timestamp 1688980957
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_204
timestamp 1688980957
transform 1 0 19872 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_219
timestamp 1688980957
transform 1 0 21252 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_235
timestamp 1688980957
transform 1 0 22724 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_247
timestamp 1688980957
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_328
timestamp 1688980957
transform 1 0 31280 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_332
timestamp 1688980957
transform 1 0 31648 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_347
timestamp 1688980957
transform 1 0 33028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_351
timestamp 1688980957
transform 1 0 33396 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_355
timestamp 1688980957
transform 1 0 33764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_369
timestamp 1688980957
transform 1 0 35052 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_381
timestamp 1688980957
transform 1 0 36156 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_392
timestamp 1688980957
transform 1 0 37168 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_400
timestamp 1688980957
transform 1 0 37904 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_23
timestamp 1688980957
transform 1 0 3220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_31
timestamp 1688980957
transform 1 0 3956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1688980957
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_63
timestamp 1688980957
transform 1 0 6900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_67
timestamp 1688980957
transform 1 0 7268 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_82
timestamp 1688980957
transform 1 0 8648 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_95
timestamp 1688980957
transform 1 0 9844 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_107
timestamp 1688980957
transform 1 0 10948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_136
timestamp 1688980957
transform 1 0 13616 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_140
timestamp 1688980957
transform 1 0 13984 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_150
timestamp 1688980957
transform 1 0 14904 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_162
timestamp 1688980957
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_190
timestamp 1688980957
transform 1 0 18584 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_253
timestamp 1688980957
transform 1 0 24380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_265
timestamp 1688980957
transform 1 0 25484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_277
timestamp 1688980957
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_296
timestamp 1688980957
transform 1 0 28336 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_302
timestamp 1688980957
transform 1 0 28888 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1688980957
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 1688980957
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 1688980957
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_345
timestamp 1688980957
transform 1 0 32844 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_368
timestamp 1688980957
transform 1 0 34960 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_376
timestamp 1688980957
transform 1 0 35696 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_380
timestamp 1688980957
transform 1 0 36064 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_10
timestamp 1688980957
transform 1 0 2024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_25
timestamp 1688980957
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 1688980957
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_102
timestamp 1688980957
transform 1 0 10488 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_110
timestamp 1688980957
transform 1 0 11224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_122
timestamp 1688980957
transform 1 0 12328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_150
timestamp 1688980957
transform 1 0 14904 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_161
timestamp 1688980957
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_216
timestamp 1688980957
transform 1 0 20976 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_228
timestamp 1688980957
transform 1 0 22080 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_256
timestamp 1688980957
transform 1 0 24656 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_282
timestamp 1688980957
transform 1 0 27048 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_294
timestamp 1688980957
transform 1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_306
timestamp 1688980957
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_316
timestamp 1688980957
transform 1 0 30176 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_340
timestamp 1688980957
transform 1 0 32384 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_348
timestamp 1688980957
transform 1 0 33120 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_354
timestamp 1688980957
transform 1 0 33672 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_362
timestamp 1688980957
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 1688980957
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_11
timestamp 1688980957
transform 1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_23
timestamp 1688980957
transform 1 0 3220 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_32
timestamp 1688980957
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_44
timestamp 1688980957
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_65
timestamp 1688980957
transform 1 0 7084 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_75
timestamp 1688980957
transform 1 0 8004 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_87
timestamp 1688980957
transform 1 0 9108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_99
timestamp 1688980957
transform 1 0 10212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_120
timestamp 1688980957
transform 1 0 12144 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_132
timestamp 1688980957
transform 1 0 13248 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_140
timestamp 1688980957
transform 1 0 13984 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_150
timestamp 1688980957
transform 1 0 14904 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_162
timestamp 1688980957
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_177
timestamp 1688980957
transform 1 0 17388 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_200
timestamp 1688980957
transform 1 0 19504 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1688980957
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_249
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_257
timestamp 1688980957
transform 1 0 24748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_264
timestamp 1688980957
transform 1 0 25392 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_275
timestamp 1688980957
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_291
timestamp 1688980957
transform 1 0 27876 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_299
timestamp 1688980957
transform 1 0 28612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_305
timestamp 1688980957
transform 1 0 29164 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_326
timestamp 1688980957
transform 1 0 31096 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_334
timestamp 1688980957
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_345
timestamp 1688980957
transform 1 0 32844 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_353
timestamp 1688980957
transform 1 0 33580 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_365
timestamp 1688980957
transform 1 0 34684 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_380
timestamp 1688980957
transform 1 0 36064 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_9
timestamp 1688980957
transform 1 0 1932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_21
timestamp 1688980957
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_36
timestamp 1688980957
transform 1 0 4416 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_44
timestamp 1688980957
transform 1 0 5152 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_50
timestamp 1688980957
transform 1 0 5704 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_62
timestamp 1688980957
transform 1 0 6808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_75
timestamp 1688980957
transform 1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_99
timestamp 1688980957
transform 1 0 10212 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_111
timestamp 1688980957
transform 1 0 11316 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_123
timestamp 1688980957
transform 1 0 12420 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_135
timestamp 1688980957
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_158
timestamp 1688980957
transform 1 0 15640 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_170
timestamp 1688980957
transform 1 0 16744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_179
timestamp 1688980957
transform 1 0 17572 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_187
timestamp 1688980957
transform 1 0 18308 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_201
timestamp 1688980957
transform 1 0 19596 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_210
timestamp 1688980957
transform 1 0 20424 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_237
timestamp 1688980957
transform 1 0 22908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_249
timestamp 1688980957
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_257
timestamp 1688980957
transform 1 0 24748 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_264
timestamp 1688980957
transform 1 0 25392 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_276
timestamp 1688980957
transform 1 0 26496 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_291
timestamp 1688980957
transform 1 0 27876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_303
timestamp 1688980957
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_315
timestamp 1688980957
transform 1 0 30084 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_322
timestamp 1688980957
transform 1 0 30728 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_334
timestamp 1688980957
transform 1 0 31832 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_346
timestamp 1688980957
transform 1 0 32936 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_358
timestamp 1688980957
transform 1 0 34040 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_376
timestamp 1688980957
transform 1 0 35696 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_388
timestamp 1688980957
transform 1 0 36800 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_40
timestamp 1688980957
transform 1 0 4784 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_80
timestamp 1688980957
transform 1 0 8464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_86
timestamp 1688980957
transform 1 0 9016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_101
timestamp 1688980957
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1688980957
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_122
timestamp 1688980957
transform 1 0 12328 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_128
timestamp 1688980957
transform 1 0 12880 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_147
timestamp 1688980957
transform 1 0 14628 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_158
timestamp 1688980957
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1688980957
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_175
timestamp 1688980957
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_190
timestamp 1688980957
transform 1 0 18584 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_210
timestamp 1688980957
transform 1 0 20424 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_222
timestamp 1688980957
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_233
timestamp 1688980957
transform 1 0 22540 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_245
timestamp 1688980957
transform 1 0 23644 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_257
timestamp 1688980957
transform 1 0 24748 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_268
timestamp 1688980957
transform 1 0 25760 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_285
timestamp 1688980957
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_290
timestamp 1688980957
transform 1 0 27784 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_302
timestamp 1688980957
transform 1 0 28888 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_310
timestamp 1688980957
transform 1 0 29624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_315
timestamp 1688980957
transform 1 0 30084 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_321
timestamp 1688980957
transform 1 0 30636 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_325
timestamp 1688980957
transform 1 0 31004 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_333
timestamp 1688980957
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_346
timestamp 1688980957
transform 1 0 32936 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_358
timestamp 1688980957
transform 1 0 34040 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_388
timestamp 1688980957
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_10
timestamp 1688980957
transform 1 0 2024 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_22
timestamp 1688980957
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_37
timestamp 1688980957
transform 1 0 4508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_49
timestamp 1688980957
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_61
timestamp 1688980957
transform 1 0 6716 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_69
timestamp 1688980957
transform 1 0 7452 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_79
timestamp 1688980957
transform 1 0 8372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_89
timestamp 1688980957
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_102
timestamp 1688980957
transform 1 0 10488 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_110
timestamp 1688980957
transform 1 0 11224 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_128
timestamp 1688980957
transform 1 0 12880 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_181
timestamp 1688980957
transform 1 0 17756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_193
timestamp 1688980957
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_213
timestamp 1688980957
transform 1 0 20700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_225
timestamp 1688980957
transform 1 0 21804 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_236
timestamp 1688980957
transform 1 0 22816 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_264
timestamp 1688980957
transform 1 0 25392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_276
timestamp 1688980957
transform 1 0 26496 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_306
timestamp 1688980957
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_331
timestamp 1688980957
transform 1 0 31556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_352
timestamp 1688980957
transform 1 0 33488 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_381
timestamp 1688980957
transform 1 0 36156 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_385
timestamp 1688980957
transform 1 0 36524 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_391
timestamp 1688980957
transform 1 0 37076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_399
timestamp 1688980957
transform 1 0 37812 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_21
timestamp 1688980957
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_33
timestamp 1688980957
transform 1 0 4140 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_41
timestamp 1688980957
transform 1 0 4876 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_62
timestamp 1688980957
transform 1 0 6808 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_70
timestamp 1688980957
transform 1 0 7544 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_78
timestamp 1688980957
transform 1 0 8280 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_90
timestamp 1688980957
transform 1 0 9384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_97
timestamp 1688980957
transform 1 0 10028 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_130
timestamp 1688980957
transform 1 0 13064 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_162
timestamp 1688980957
transform 1 0 16008 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_185
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_197
timestamp 1688980957
transform 1 0 19228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_215
timestamp 1688980957
transform 1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_255
timestamp 1688980957
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_263
timestamp 1688980957
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_269
timestamp 1688980957
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_277
timestamp 1688980957
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_294
timestamp 1688980957
transform 1 0 28152 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_306
timestamp 1688980957
transform 1 0 29256 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_322
timestamp 1688980957
transform 1 0 30728 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_334
timestamp 1688980957
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_340
timestamp 1688980957
transform 1 0 32384 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_355
timestamp 1688980957
transform 1 0 33764 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_367
timestamp 1688980957
transform 1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_374
timestamp 1688980957
transform 1 0 35512 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1688980957
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_396
timestamp 1688980957
transform 1 0 37536 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_10
timestamp 1688980957
transform 1 0 2024 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_33
timestamp 1688980957
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_96
timestamp 1688980957
transform 1 0 9936 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_128
timestamp 1688980957
transform 1 0 12880 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_146
timestamp 1688980957
transform 1 0 14536 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_162
timestamp 1688980957
transform 1 0 16008 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1688980957
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_215
timestamp 1688980957
transform 1 0 20884 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_229
timestamp 1688980957
transform 1 0 22172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_249
timestamp 1688980957
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_266
timestamp 1688980957
transform 1 0 25576 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_274
timestamp 1688980957
transform 1 0 26312 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_286
timestamp 1688980957
transform 1 0 27416 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_298
timestamp 1688980957
transform 1 0 28520 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1688980957
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_315
timestamp 1688980957
transform 1 0 30084 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_327
timestamp 1688980957
transform 1 0 31188 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_350
timestamp 1688980957
transform 1 0 33304 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_362
timestamp 1688980957
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_384
timestamp 1688980957
transform 1 0 36432 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_396
timestamp 1688980957
transform 1 0 37536 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_400
timestamp 1688980957
transform 1 0 37904 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_50
timestamp 1688980957
transform 1 0 5704 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_66
timestamp 1688980957
transform 1 0 7176 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_78
timestamp 1688980957
transform 1 0 8280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_131
timestamp 1688980957
transform 1 0 13156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_157
timestamp 1688980957
transform 1 0 15548 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_163
timestamp 1688980957
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_173
timestamp 1688980957
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_190
timestamp 1688980957
transform 1 0 18584 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_209
timestamp 1688980957
transform 1 0 20332 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_213
timestamp 1688980957
transform 1 0 20700 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_220
timestamp 1688980957
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_248
timestamp 1688980957
transform 1 0 23920 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_274
timestamp 1688980957
transform 1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_340
timestamp 1688980957
transform 1 0 32384 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_351
timestamp 1688980957
transform 1 0 33396 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_363
timestamp 1688980957
transform 1 0 34500 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_380
timestamp 1688980957
transform 1 0 36064 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_393
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_10
timestamp 1688980957
transform 1 0 2024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_22
timestamp 1688980957
transform 1 0 3128 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_38
timestamp 1688980957
transform 1 0 4600 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_44
timestamp 1688980957
transform 1 0 5152 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_73
timestamp 1688980957
transform 1 0 7820 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_88
timestamp 1688980957
transform 1 0 9200 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_100
timestamp 1688980957
transform 1 0 10304 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_112
timestamp 1688980957
transform 1 0 11408 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_124
timestamp 1688980957
transform 1 0 12512 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_130
timestamp 1688980957
transform 1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_134
timestamp 1688980957
transform 1 0 13432 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_155
timestamp 1688980957
transform 1 0 15364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_167
timestamp 1688980957
transform 1 0 16468 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_179
timestamp 1688980957
transform 1 0 17572 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_215
timestamp 1688980957
transform 1 0 20884 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_264
timestamp 1688980957
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_287
timestamp 1688980957
transform 1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_291
timestamp 1688980957
transform 1 0 27876 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1688980957
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_317
timestamp 1688980957
transform 1 0 30268 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_341
timestamp 1688980957
transform 1 0 32476 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 1688980957
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 1688980957
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_24
timestamp 1688980957
transform 1 0 3312 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_32
timestamp 1688980957
transform 1 0 4048 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_44
timestamp 1688980957
transform 1 0 5152 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1688980957
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_65
timestamp 1688980957
transform 1 0 7084 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_97
timestamp 1688980957
transform 1 0 10028 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_102
timestamp 1688980957
transform 1 0 10488 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_106
timestamp 1688980957
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_119
timestamp 1688980957
transform 1 0 12052 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_132
timestamp 1688980957
transform 1 0 13248 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_140
timestamp 1688980957
transform 1 0 13984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_166
timestamp 1688980957
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_183
timestamp 1688980957
transform 1 0 17940 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_254
timestamp 1688980957
transform 1 0 24472 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_266
timestamp 1688980957
transform 1 0 25576 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_290
timestamp 1688980957
transform 1 0 27784 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_298
timestamp 1688980957
transform 1 0 28520 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_325
timestamp 1688980957
transform 1 0 31004 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_345
timestamp 1688980957
transform 1 0 32844 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_353
timestamp 1688980957
transform 1 0 33580 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_359
timestamp 1688980957
transform 1 0 34132 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_369
timestamp 1688980957
transform 1 0 35052 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_381
timestamp 1688980957
transform 1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_389
timestamp 1688980957
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_7
timestamp 1688980957
transform 1 0 1748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_33
timestamp 1688980957
transform 1 0 4140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_45
timestamp 1688980957
transform 1 0 5244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_57
timestamp 1688980957
transform 1 0 6348 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_71
timestamp 1688980957
transform 1 0 7636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_135
timestamp 1688980957
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_145
timestamp 1688980957
transform 1 0 14444 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_152
timestamp 1688980957
transform 1 0 15088 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_160
timestamp 1688980957
transform 1 0 15824 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_178
timestamp 1688980957
transform 1 0 17480 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_186
timestamp 1688980957
transform 1 0 18216 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_225
timestamp 1688980957
transform 1 0 21804 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_237
timestamp 1688980957
transform 1 0 22908 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_250
timestamp 1688980957
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_264
timestamp 1688980957
transform 1 0 25392 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_276
timestamp 1688980957
transform 1 0 26496 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_282
timestamp 1688980957
transform 1 0 27048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_291
timestamp 1688980957
transform 1 0 27876 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_306
timestamp 1688980957
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_313
timestamp 1688980957
transform 1 0 29900 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_322
timestamp 1688980957
transform 1 0 30728 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_334
timestamp 1688980957
transform 1 0 31832 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_346
timestamp 1688980957
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_358
timestamp 1688980957
transform 1 0 34040 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_388
timestamp 1688980957
transform 1 0 36800 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_400
timestamp 1688980957
transform 1 0 37904 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_9
timestamp 1688980957
transform 1 0 1932 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_17
timestamp 1688980957
transform 1 0 2668 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_22
timestamp 1688980957
transform 1 0 3128 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_44
timestamp 1688980957
transform 1 0 5152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_50
timestamp 1688980957
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_103
timestamp 1688980957
transform 1 0 10580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_204
timestamp 1688980957
transform 1 0 19872 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_229
timestamp 1688980957
transform 1 0 22172 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_253
timestamp 1688980957
transform 1 0 24380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_278
timestamp 1688980957
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1688980957
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_354
timestamp 1688980957
transform 1 0 33672 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 1688980957
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 1688980957
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1688980957
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_88
timestamp 1688980957
transform 1 0 9200 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_100
timestamp 1688980957
transform 1 0 10304 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_112
timestamp 1688980957
transform 1 0 11408 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_124
timestamp 1688980957
transform 1 0 12512 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_159
timestamp 1688980957
transform 1 0 15732 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_167
timestamp 1688980957
transform 1 0 16468 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_178
timestamp 1688980957
transform 1 0 17480 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_190
timestamp 1688980957
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_205
timestamp 1688980957
transform 1 0 19964 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_213
timestamp 1688980957
transform 1 0 20700 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_241
timestamp 1688980957
transform 1 0 23276 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_248
timestamp 1688980957
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_261
timestamp 1688980957
transform 1 0 25116 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_278
timestamp 1688980957
transform 1 0 26680 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_299
timestamp 1688980957
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_318
timestamp 1688980957
transform 1 0 30360 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_348
timestamp 1688980957
transform 1 0 33120 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_358
timestamp 1688980957
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_391
timestamp 1688980957
transform 1 0 37076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_399
timestamp 1688980957
transform 1 0 37812 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_102
timestamp 1688980957
transform 1 0 10488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_110
timestamp 1688980957
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_129
timestamp 1688980957
transform 1 0 12972 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_141
timestamp 1688980957
transform 1 0 14076 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_151
timestamp 1688980957
transform 1 0 14996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_155
timestamp 1688980957
transform 1 0 15364 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_160
timestamp 1688980957
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_176
timestamp 1688980957
transform 1 0 17296 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_185
timestamp 1688980957
transform 1 0 18124 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_191
timestamp 1688980957
transform 1 0 18676 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_197
timestamp 1688980957
transform 1 0 19228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_209
timestamp 1688980957
transform 1 0 20332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_221
timestamp 1688980957
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_236
timestamp 1688980957
transform 1 0 22816 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_248
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_260
timestamp 1688980957
transform 1 0 25024 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_268
timestamp 1688980957
transform 1 0 25760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_284
timestamp 1688980957
transform 1 0 27232 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_333
timestamp 1688980957
transform 1 0 31740 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_345
timestamp 1688980957
transform 1 0 32844 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_374
timestamp 1688980957
transform 1 0 35512 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_386
timestamp 1688980957
transform 1 0 36616 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_37
timestamp 1688980957
transform 1 0 4508 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_64
timestamp 1688980957
transform 1 0 6992 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_76
timestamp 1688980957
transform 1 0 8096 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_123
timestamp 1688980957
transform 1 0 12420 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_148
timestamp 1688980957
transform 1 0 14720 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_156
timestamp 1688980957
transform 1 0 15456 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_163
timestamp 1688980957
transform 1 0 16100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_194
timestamp 1688980957
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_233
timestamp 1688980957
transform 1 0 22540 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_247
timestamp 1688980957
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_295
timestamp 1688980957
transform 1 0 28244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1688980957
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_315
timestamp 1688980957
transform 1 0 30084 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_326
timestamp 1688980957
transform 1 0 31096 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_338
timestamp 1688980957
transform 1 0 32200 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_350
timestamp 1688980957
transform 1 0 33304 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_358
timestamp 1688980957
transform 1 0 34040 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1688980957
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_31
timestamp 1688980957
transform 1 0 3956 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_53
timestamp 1688980957
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_66
timestamp 1688980957
transform 1 0 7176 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_70
timestamp 1688980957
transform 1 0 7544 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_101
timestamp 1688980957
transform 1 0 10396 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_106
timestamp 1688980957
transform 1 0 10856 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_122
timestamp 1688980957
transform 1 0 12328 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_130
timestamp 1688980957
transform 1 0 13064 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_134
timestamp 1688980957
transform 1 0 13432 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_151
timestamp 1688980957
transform 1 0 14996 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_163
timestamp 1688980957
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_177
timestamp 1688980957
transform 1 0 17388 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_189
timestamp 1688980957
transform 1 0 18492 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1688980957
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_255
timestamp 1688980957
transform 1 0 24564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_267
timestamp 1688980957
transform 1 0 25668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_347
timestamp 1688980957
transform 1 0 33028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_359
timestamp 1688980957
transform 1 0 34132 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_363
timestamp 1688980957
transform 1 0 34500 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_369
timestamp 1688980957
transform 1 0 35052 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_381
timestamp 1688980957
transform 1 0 36156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_389
timestamp 1688980957
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_397
timestamp 1688980957
transform 1 0 37628 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_36
timestamp 1688980957
transform 1 0 4416 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_40
timestamp 1688980957
transform 1 0 4784 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_79
timestamp 1688980957
transform 1 0 8372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_93
timestamp 1688980957
transform 1 0 9660 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_119
timestamp 1688980957
transform 1 0 12052 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_131
timestamp 1688980957
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_161
timestamp 1688980957
transform 1 0 15916 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_170
timestamp 1688980957
transform 1 0 16744 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_182
timestamp 1688980957
transform 1 0 17848 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_194
timestamp 1688980957
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_207
timestamp 1688980957
transform 1 0 20148 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_213
timestamp 1688980957
transform 1 0 20700 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_234
timestamp 1688980957
transform 1 0 22632 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_246
timestamp 1688980957
transform 1 0 23736 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_260
timestamp 1688980957
transform 1 0 25024 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_275
timestamp 1688980957
transform 1 0 26404 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_287
timestamp 1688980957
transform 1 0 27508 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_299
timestamp 1688980957
transform 1 0 28612 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_303
timestamp 1688980957
transform 1 0 28980 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_332
timestamp 1688980957
transform 1 0 31648 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_354
timestamp 1688980957
transform 1 0 33672 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_386
timestamp 1688980957
transform 1 0 36616 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_398
timestamp 1688980957
transform 1 0 37720 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_53
timestamp 1688980957
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_68
timestamp 1688980957
transform 1 0 7360 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_79
timestamp 1688980957
transform 1 0 8372 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_133
timestamp 1688980957
transform 1 0 13340 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_145
timestamp 1688980957
transform 1 0 14444 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_157
timestamp 1688980957
transform 1 0 15548 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_165
timestamp 1688980957
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_194
timestamp 1688980957
transform 1 0 18952 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_206
timestamp 1688980957
transform 1 0 20056 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_212
timestamp 1688980957
transform 1 0 20608 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_220
timestamp 1688980957
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_241
timestamp 1688980957
transform 1 0 23276 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_250
timestamp 1688980957
transform 1 0 24104 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_262
timestamp 1688980957
transform 1 0 25208 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_326
timestamp 1688980957
transform 1 0 31096 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_348
timestamp 1688980957
transform 1 0 33120 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_360
timestamp 1688980957
transform 1 0 34224 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_370
timestamp 1688980957
transform 1 0 35144 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_382
timestamp 1688980957
transform 1 0 36248 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 1688980957
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_34
timestamp 1688980957
transform 1 0 4232 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_46
timestamp 1688980957
transform 1 0 5336 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_56
timestamp 1688980957
transform 1 0 6256 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_68
timestamp 1688980957
transform 1 0 7360 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_76
timestamp 1688980957
transform 1 0 8096 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_106
timestamp 1688980957
transform 1 0 10856 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_118
timestamp 1688980957
transform 1 0 11960 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_129
timestamp 1688980957
transform 1 0 12972 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_149
timestamp 1688980957
transform 1 0 14812 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_166
timestamp 1688980957
transform 1 0 16376 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_176
timestamp 1688980957
transform 1 0 17296 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_184
timestamp 1688980957
transform 1 0 18032 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_194
timestamp 1688980957
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_219
timestamp 1688980957
transform 1 0 21252 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_231
timestamp 1688980957
transform 1 0 22356 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_243
timestamp 1688980957
transform 1 0 23460 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_250
timestamp 1688980957
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_258
timestamp 1688980957
transform 1 0 24840 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_264
timestamp 1688980957
transform 1 0 25392 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_280
timestamp 1688980957
transform 1 0 26864 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_299
timestamp 1688980957
transform 1 0 28612 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_325
timestamp 1688980957
transform 1 0 31004 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_347
timestamp 1688980957
transform 1 0 33028 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 1688980957
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_33
timestamp 1688980957
transform 1 0 4140 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_76
timestamp 1688980957
transform 1 0 8096 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_80
timestamp 1688980957
transform 1 0 8464 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_84
timestamp 1688980957
transform 1 0 8832 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_96
timestamp 1688980957
transform 1 0 9936 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_108
timestamp 1688980957
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_122
timestamp 1688980957
transform 1 0 12328 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_128
timestamp 1688980957
transform 1 0 12880 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_177
timestamp 1688980957
transform 1 0 17388 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_201
timestamp 1688980957
transform 1 0 19596 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_216
timestamp 1688980957
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_241
timestamp 1688980957
transform 1 0 23276 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_262
timestamp 1688980957
transform 1 0 25208 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_266
timestamp 1688980957
transform 1 0 25576 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_274
timestamp 1688980957
transform 1 0 26312 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_319
timestamp 1688980957
transform 1 0 30452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_331
timestamp 1688980957
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_345
timestamp 1688980957
transform 1 0 32844 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_357
timestamp 1688980957
transform 1 0 33948 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_369
timestamp 1688980957
transform 1 0 35052 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_381
timestamp 1688980957
transform 1 0 36156 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_389
timestamp 1688980957
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_38
timestamp 1688980957
transform 1 0 4600 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_46
timestamp 1688980957
transform 1 0 5336 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_82
timestamp 1688980957
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_94
timestamp 1688980957
transform 1 0 9752 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_106
timestamp 1688980957
transform 1 0 10856 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_118
timestamp 1688980957
transform 1 0 11960 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_130
timestamp 1688980957
transform 1 0 13064 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_150
timestamp 1688980957
transform 1 0 14904 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_162
timestamp 1688980957
transform 1 0 16008 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_225
timestamp 1688980957
transform 1 0 21804 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_237
timestamp 1688980957
transform 1 0 22908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_249
timestamp 1688980957
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_259
timestamp 1688980957
transform 1 0 24932 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_278
timestamp 1688980957
transform 1 0 26680 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_290
timestamp 1688980957
transform 1 0 27784 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_302
timestamp 1688980957
transform 1 0 28888 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_344
timestamp 1688980957
transform 1 0 32752 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_359
timestamp 1688980957
transform 1 0 34132 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_374
timestamp 1688980957
transform 1 0 35512 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_386
timestamp 1688980957
transform 1 0 36616 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_398
timestamp 1688980957
transform 1 0 37720 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_94
timestamp 1688980957
transform 1 0 9752 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_107
timestamp 1688980957
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_120
timestamp 1688980957
transform 1 0 12144 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_128
timestamp 1688980957
transform 1 0 12880 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_184
timestamp 1688980957
transform 1 0 18032 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_206
timestamp 1688980957
transform 1 0 20056 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_232
timestamp 1688980957
transform 1 0 22448 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_386
timestamp 1688980957
transform 1 0 36616 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_57
timestamp 1688980957
transform 1 0 6348 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_81
timestamp 1688980957
transform 1 0 8556 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_111
timestamp 1688980957
transform 1 0 11316 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_123
timestamp 1688980957
transform 1 0 12420 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_129
timestamp 1688980957
transform 1 0 12972 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_137
timestamp 1688980957
transform 1 0 13708 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_220
timestamp 1688980957
transform 1 0 21344 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_250
timestamp 1688980957
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_267
timestamp 1688980957
transform 1 0 25668 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_282
timestamp 1688980957
transform 1 0 27048 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_296
timestamp 1688980957
transform 1 0 28336 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_320
timestamp 1688980957
transform 1 0 30544 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_328
timestamp 1688980957
transform 1 0 31280 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_336
timestamp 1688980957
transform 1 0 32016 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_348
timestamp 1688980957
transform 1 0 33120 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_360
timestamp 1688980957
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_374
timestamp 1688980957
transform 1 0 35512 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_386
timestamp 1688980957
transform 1 0 36616 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_398
timestamp 1688980957
transform 1 0 37720 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_45
timestamp 1688980957
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_53
timestamp 1688980957
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_120
timestamp 1688980957
transform 1 0 12144 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_126
timestamp 1688980957
transform 1 0 12696 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_138
timestamp 1688980957
transform 1 0 13800 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_150
timestamp 1688980957
transform 1 0 14904 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_162
timestamp 1688980957
transform 1 0 16008 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_175
timestamp 1688980957
transform 1 0 17204 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_182
timestamp 1688980957
transform 1 0 17848 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_186
timestamp 1688980957
transform 1 0 18216 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_195
timestamp 1688980957
transform 1 0 19044 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_199
timestamp 1688980957
transform 1 0 19412 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_220
timestamp 1688980957
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_231
timestamp 1688980957
transform 1 0 22356 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_235
timestamp 1688980957
transform 1 0 22724 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_243
timestamp 1688980957
transform 1 0 23460 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_253
timestamp 1688980957
transform 1 0 24380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_265
timestamp 1688980957
transform 1 0 25484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_277
timestamp 1688980957
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_292
timestamp 1688980957
transform 1 0 27968 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_306
timestamp 1688980957
transform 1 0 29256 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_318
timestamp 1688980957
transform 1 0 30360 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_331
timestamp 1688980957
transform 1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_354
timestamp 1688980957
transform 1 0 33672 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_366
timestamp 1688980957
transform 1 0 34776 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_374
timestamp 1688980957
transform 1 0 35512 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_380
timestamp 1688980957
transform 1 0 36064 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_81
timestamp 1688980957
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_89
timestamp 1688980957
transform 1 0 9292 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_99
timestamp 1688980957
transform 1 0 10212 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_111
timestamp 1688980957
transform 1 0 11316 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_123
timestamp 1688980957
transform 1 0 12420 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_135
timestamp 1688980957
transform 1 0 13524 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_161
timestamp 1688980957
transform 1 0 15916 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_179
timestamp 1688980957
transform 1 0 17572 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_193
timestamp 1688980957
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_205
timestamp 1688980957
transform 1 0 19964 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_214
timestamp 1688980957
transform 1 0 20792 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_231
timestamp 1688980957
transform 1 0 22356 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_239
timestamp 1688980957
transform 1 0 23092 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_286
timestamp 1688980957
transform 1 0 27416 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_315
timestamp 1688980957
transform 1 0 30084 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_319
timestamp 1688980957
transform 1 0 30452 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_323
timestamp 1688980957
transform 1 0 30820 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_348
timestamp 1688980957
transform 1 0 33120 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_360
timestamp 1688980957
transform 1 0 34224 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_388
timestamp 1688980957
transform 1 0 36800 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_400
timestamp 1688980957
transform 1 0 37904 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_63
timestamp 1688980957
transform 1 0 6900 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_106
timestamp 1688980957
transform 1 0 10856 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_147
timestamp 1688980957
transform 1 0 14628 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_159
timestamp 1688980957
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_180
timestamp 1688980957
transform 1 0 17664 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_192
timestamp 1688980957
transform 1 0 18768 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_222
timestamp 1688980957
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_228
timestamp 1688980957
transform 1 0 22080 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_240
timestamp 1688980957
transform 1 0 23184 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_251
timestamp 1688980957
transform 1 0 24196 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_257
timestamp 1688980957
transform 1 0 24748 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_265
timestamp 1688980957
transform 1 0 25484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_304
timestamp 1688980957
transform 1 0 29072 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_316
timestamp 1688980957
transform 1 0 30176 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_328
timestamp 1688980957
transform 1 0 31280 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_345
timestamp 1688980957
transform 1 0 32844 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_368
timestamp 1688980957
transform 1 0 34960 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_380
timestamp 1688980957
transform 1 0 36064 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_386
timestamp 1688980957
transform 1 0 36616 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_390
timestamp 1688980957
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_37
timestamp 1688980957
transform 1 0 4508 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_63
timestamp 1688980957
transform 1 0 6900 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_68
timestamp 1688980957
transform 1 0 7360 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_80
timestamp 1688980957
transform 1 0 8464 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_96
timestamp 1688980957
transform 1 0 9936 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_108
timestamp 1688980957
transform 1 0 11040 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_118
timestamp 1688980957
transform 1 0 11960 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_130
timestamp 1688980957
transform 1 0 13064 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_138
timestamp 1688980957
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_170
timestamp 1688980957
transform 1 0 16744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_178
timestamp 1688980957
transform 1 0 17480 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_201
timestamp 1688980957
transform 1 0 19596 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_211
timestamp 1688980957
transform 1 0 20516 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_229
timestamp 1688980957
transform 1 0 22172 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_248
timestamp 1688980957
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_261
timestamp 1688980957
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_278
timestamp 1688980957
transform 1 0 26680 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_285
timestamp 1688980957
transform 1 0 27324 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_294
timestamp 1688980957
transform 1 0 28152 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_306
timestamp 1688980957
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_317
timestamp 1688980957
transform 1 0 30268 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_327
timestamp 1688980957
transform 1 0 31188 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_336
timestamp 1688980957
transform 1 0 32016 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_348
timestamp 1688980957
transform 1 0 33120 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_359
timestamp 1688980957
transform 1 0 34132 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_388
timestamp 1688980957
transform 1 0 36800 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_400
timestamp 1688980957
transform 1 0 37904 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_50
timestamp 1688980957
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_83
timestamp 1688980957
transform 1 0 8740 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_95
timestamp 1688980957
transform 1 0 9844 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_107
timestamp 1688980957
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_121
timestamp 1688980957
transform 1 0 12236 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_133
timestamp 1688980957
transform 1 0 13340 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_145
timestamp 1688980957
transform 1 0 14444 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_157
timestamp 1688980957
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_165
timestamp 1688980957
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_177
timestamp 1688980957
transform 1 0 17388 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_189
timestamp 1688980957
transform 1 0 18492 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_201
timestamp 1688980957
transform 1 0 19596 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_213
timestamp 1688980957
transform 1 0 20700 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_221
timestamp 1688980957
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_234
timestamp 1688980957
transform 1 0 22632 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_320
timestamp 1688980957
transform 1 0 30544 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_326
timestamp 1688980957
transform 1 0 31096 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_345
timestamp 1688980957
transform 1 0 32844 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_355
timestamp 1688980957
transform 1 0 33764 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_367
timestamp 1688980957
transform 1 0 34868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_379
timestamp 1688980957
transform 1 0 35972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1688980957
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_59
timestamp 1688980957
transform 1 0 6532 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_100
timestamp 1688980957
transform 1 0 10304 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_112
timestamp 1688980957
transform 1 0 11408 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_124
timestamp 1688980957
transform 1 0 12512 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_136
timestamp 1688980957
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_173
timestamp 1688980957
transform 1 0 17020 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_179
timestamp 1688980957
transform 1 0 17572 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_191
timestamp 1688980957
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_249
timestamp 1688980957
transform 1 0 24012 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_261
timestamp 1688980957
transform 1 0 25116 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_279
timestamp 1688980957
transform 1 0 26772 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_297
timestamp 1688980957
transform 1 0 28428 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_303
timestamp 1688980957
transform 1 0 28980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_317
timestamp 1688980957
transform 1 0 30268 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_342
timestamp 1688980957
transform 1 0 32568 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1688980957
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1688980957
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_62
timestamp 1688980957
transform 1 0 6808 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_66
timestamp 1688980957
transform 1 0 7176 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_109
timestamp 1688980957
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_151
timestamp 1688980957
transform 1 0 14996 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_163
timestamp 1688980957
transform 1 0 16100 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_189
timestamp 1688980957
transform 1 0 18492 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_199
timestamp 1688980957
transform 1 0 19412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_211
timestamp 1688980957
transform 1 0 20516 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_221
timestamp 1688980957
transform 1 0 21436 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_234
timestamp 1688980957
transform 1 0 22632 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_251
timestamp 1688980957
transform 1 0 24196 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_257
timestamp 1688980957
transform 1 0 24748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_285
timestamp 1688980957
transform 1 0 27324 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_307
timestamp 1688980957
transform 1 0 29348 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_324
timestamp 1688980957
transform 1 0 30912 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_330
timestamp 1688980957
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_343
timestamp 1688980957
transform 1 0 32660 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_347
timestamp 1688980957
transform 1 0 33028 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_353
timestamp 1688980957
transform 1 0 33580 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_365
timestamp 1688980957
transform 1 0 34684 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_377
timestamp 1688980957
transform 1 0 35788 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_389
timestamp 1688980957
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_49
timestamp 1688980957
transform 1 0 5612 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_74
timestamp 1688980957
transform 1 0 7912 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_82
timestamp 1688980957
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_95
timestamp 1688980957
transform 1 0 9844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_107
timestamp 1688980957
transform 1 0 10948 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_134
timestamp 1688980957
transform 1 0 13432 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_150
timestamp 1688980957
transform 1 0 14904 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_168
timestamp 1688980957
transform 1 0 16560 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_185
timestamp 1688980957
transform 1 0 18124 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_192
timestamp 1688980957
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_233
timestamp 1688980957
transform 1 0 22540 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_241
timestamp 1688980957
transform 1 0 23276 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1688980957
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_272
timestamp 1688980957
transform 1 0 26128 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_292
timestamp 1688980957
transform 1 0 27968 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_339
timestamp 1688980957
transform 1 0 32292 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_351
timestamp 1688980957
transform 1 0 33396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1688980957
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_65
timestamp 1688980957
transform 1 0 7084 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_72
timestamp 1688980957
transform 1 0 7728 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_84
timestamp 1688980957
transform 1 0 8832 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_88
timestamp 1688980957
transform 1 0 9200 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_98
timestamp 1688980957
transform 1 0 10120 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_110
timestamp 1688980957
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_205
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_213
timestamp 1688980957
transform 1 0 20700 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_218
timestamp 1688980957
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_237
timestamp 1688980957
transform 1 0 22908 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_250
timestamp 1688980957
transform 1 0 24104 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_260
timestamp 1688980957
transform 1 0 25024 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_272
timestamp 1688980957
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_290
timestamp 1688980957
transform 1 0 27784 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_298
timestamp 1688980957
transform 1 0 28520 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_304
timestamp 1688980957
transform 1 0 29072 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_314
timestamp 1688980957
transform 1 0 29992 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1688980957
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_360
timestamp 1688980957
transform 1 0 34224 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_372
timestamp 1688980957
transform 1 0 35328 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_384
timestamp 1688980957
transform 1 0 36432 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_7
timestamp 1688980957
transform 1 0 1748 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_19
timestamp 1688980957
transform 1 0 2852 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_106
timestamp 1688980957
transform 1 0 10856 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_118
timestamp 1688980957
transform 1 0 11960 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_130
timestamp 1688980957
transform 1 0 13064 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_138
timestamp 1688980957
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_177
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_192
timestamp 1688980957
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_205
timestamp 1688980957
transform 1 0 19964 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_240
timestamp 1688980957
transform 1 0 23184 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_248
timestamp 1688980957
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_265
timestamp 1688980957
transform 1 0 25484 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_280
timestamp 1688980957
transform 1 0 26864 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_284
timestamp 1688980957
transform 1 0 27232 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_294
timestamp 1688980957
transform 1 0 28152 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_306
timestamp 1688980957
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_334
timestamp 1688980957
transform 1 0 31832 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_343
timestamp 1688980957
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_355
timestamp 1688980957
transform 1 0 33764 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1688980957
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_97
timestamp 1688980957
transform 1 0 10028 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_108
timestamp 1688980957
transform 1 0 11040 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_131
timestamp 1688980957
transform 1 0 13156 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1688980957
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_174
timestamp 1688980957
transform 1 0 17112 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_182
timestamp 1688980957
transform 1 0 17848 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_194
timestamp 1688980957
transform 1 0 18952 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_198
timestamp 1688980957
transform 1 0 19320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1688980957
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_236
timestamp 1688980957
transform 1 0 22816 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_254
timestamp 1688980957
transform 1 0 24472 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_276
timestamp 1688980957
transform 1 0 26496 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_281
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_297
timestamp 1688980957
transform 1 0 28428 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_328
timestamp 1688980957
transform 1 0 31280 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1688980957
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 1688980957
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 1688980957
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 1688980957
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 1688980957
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_393
timestamp 1688980957
transform 1 0 37260 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_45
timestamp 1688980957
transform 1 0 5244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_57
timestamp 1688980957
transform 1 0 6348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_69
timestamp 1688980957
transform 1 0 7452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_110
timestamp 1688980957
transform 1 0 11224 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_134
timestamp 1688980957
transform 1 0 13432 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_185
timestamp 1688980957
transform 1 0 18124 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_190
timestamp 1688980957
transform 1 0 18584 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_217
timestamp 1688980957
transform 1 0 21068 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 1688980957
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_259
timestamp 1688980957
transform 1 0 24932 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 1688980957
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_312
timestamp 1688980957
transform 1 0 29808 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_324
timestamp 1688980957
transform 1 0 30912 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_339
timestamp 1688980957
transform 1 0 32292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_351
timestamp 1688980957
transform 1 0 33396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1688980957
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_368
timestamp 1688980957
transform 1 0 34960 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_380
timestamp 1688980957
transform 1 0 36064 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_392
timestamp 1688980957
transform 1 0 37168 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_9
timestamp 1688980957
transform 1 0 1932 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_21
timestamp 1688980957
transform 1 0 3036 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_29
timestamp 1688980957
transform 1 0 3772 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_37
timestamp 1688980957
transform 1 0 4508 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_44
timestamp 1688980957
transform 1 0 5152 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_85
timestamp 1688980957
transform 1 0 8924 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_122
timestamp 1688980957
transform 1 0 12328 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_128
timestamp 1688980957
transform 1 0 12880 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_133
timestamp 1688980957
transform 1 0 13340 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_139
timestamp 1688980957
transform 1 0 13892 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_141
timestamp 1688980957
transform 1 0 14076 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_153
timestamp 1688980957
transform 1 0 15180 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_177
timestamp 1688980957
transform 1 0 17388 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_184
timestamp 1688980957
transform 1 0 18032 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_197
timestamp 1688980957
transform 1 0 19228 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_202
timestamp 1688980957
transform 1 0 19688 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_216
timestamp 1688980957
transform 1 0 20976 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_233
timestamp 1688980957
transform 1 0 22540 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_245
timestamp 1688980957
transform 1 0 23644 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_251
timestamp 1688980957
transform 1 0 24196 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_253
timestamp 1688980957
transform 1 0 24380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_265
timestamp 1688980957
transform 1 0 25484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_277
timestamp 1688980957
transform 1 0 26588 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_290
timestamp 1688980957
transform 1 0 27784 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_302
timestamp 1688980957
transform 1 0 28888 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_309
timestamp 1688980957
transform 1 0 29532 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_321
timestamp 1688980957
transform 1 0 30636 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 1688980957
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 1688980957
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_337
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_345
timestamp 1688980957
transform 1 0 32844 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_352
timestamp 1688980957
transform 1 0 33488 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_365
timestamp 1688980957
transform 1 0 34684 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_373
timestamp 1688980957
transform 1 0 35420 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_380
timestamp 1688980957
transform 1 0 36064 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_393
timestamp 1688980957
transform 1 0 37260 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_399
timestamp 1688980957
transform 1 0 37812 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 9476 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 13524 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 15272 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 9660 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 8372 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 6716 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 6532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 11316 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 12696 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1688980957
transform -1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1688980957
transform -1 0 31372 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1688980957
transform -1 0 11408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1688980957
transform -1 0 15916 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1688980957
transform 1 0 37444 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1688980957
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  max_cap47
timestamp 1688980957
transform -1 0 6256 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap48
timestamp 1688980957
transform -1 0 23460 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  max_cap49
timestamp 1688980957
transform 1 0 22816 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  max_cap52
timestamp 1688980957
transform 1 0 17112 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  max_cap53
timestamp 1688980957
transform 1 0 14536 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap54
timestamp 1688980957
transform -1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  max_cap55
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  max_cap56
timestamp 1688980957
transform 1 0 15916 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1688980957
transform -1 0 18032 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1688980957
transform -1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1688980957
transform 1 0 37444 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1688980957
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1688980957
transform 1 0 37628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1688980957
transform -1 0 1932 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1688980957
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform -1 0 1932 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform -1 0 22540 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform -1 0 1932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform 1 0 37444 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1688980957
transform 1 0 12972 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform -1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform -1 0 2576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1688980957
transform 1 0 37628 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform -1 0 1932 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 37444 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 37444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1688980957
transform 1 0 9108 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform 1 0 37444 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform -1 0 7084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform -1 0 1932 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1688980957
transform 1 0 37628 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform -1 0 19964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 35512 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform 1 0 32936 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1688980957
transform -1 0 5152 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1688980957
transform -1 0 12052 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output44
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output45
timestamp 1688980957
transform -1 0 1932 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output46
timestamp 1688980957
transform 1 0 37444 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 38272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 38272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 38272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 38272 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 38272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 38272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 38272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 38272 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 38272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 38272 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 38272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 38272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 38272 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 38272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 38272 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 38272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 38272 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 38272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 38272 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 38272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 38272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 38272 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 38272 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 38272 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 38272 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 38272 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 38272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 38272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 38272 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 38272 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 38272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 38272 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 38272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 38272 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 38272 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 38272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 38272 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 38272 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 38272 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 38272 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 38272 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 38272 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 38272 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 38272 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 38272 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 38272 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 38272 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 38272 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 38272 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 38272 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 38272 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 38272 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 38272 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 38272 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 38272 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 38272 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 38272 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 38272 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 38272 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 38272 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 38272 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 38272 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 38272 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 38272 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 38272 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 38272 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 38272 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 38272 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 3680 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 8832 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 13984 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 19136 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 24288 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 29440 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 34592 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire50
timestamp 1688980957
transform -1 0 17572 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  wire51
timestamp 1688980957
transform -1 0 15824 0 -1 27200
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 38618 8848 39418 8968 0 FreeSans 480 0 0 0 cs
port 1 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 gpi[0]
port 2 nsew signal input
flabel metal3 s 38618 29248 39418 29368 0 FreeSans 480 0 0 0 gpi[10]
port 3 nsew signal input
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 gpi[11]
port 4 nsew signal input
flabel metal3 s 38618 13608 39418 13728 0 FreeSans 480 0 0 0 gpi[12]
port 5 nsew signal input
flabel metal2 s 1950 40762 2006 41562 0 FreeSans 224 90 0 0 gpi[13]
port 6 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 gpi[14]
port 7 nsew signal input
flabel metal3 s 38618 25168 39418 25288 0 FreeSans 480 0 0 0 gpi[15]
port 8 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 gpi[16]
port 9 nsew signal input
flabel metal3 s 38618 4088 39418 4208 0 FreeSans 480 0 0 0 gpi[17]
port 10 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 gpi[18]
port 11 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 gpi[19]
port 12 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 gpi[1]
port 13 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 gpi[20]
port 14 nsew signal input
flabel metal3 s 38618 6128 39418 6248 0 FreeSans 480 0 0 0 gpi[21]
port 15 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 gpi[22]
port 16 nsew signal input
flabel metal2 s 30930 40762 30986 41562 0 FreeSans 224 90 0 0 gpi[23]
port 17 nsew signal input
flabel metal2 s 28354 40762 28410 41562 0 FreeSans 224 90 0 0 gpi[24]
port 18 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 gpi[25]
port 19 nsew signal input
flabel metal3 s 38618 27208 39418 27328 0 FreeSans 480 0 0 0 gpi[26]
port 20 nsew signal input
flabel metal3 s 38618 31968 39418 32088 0 FreeSans 480 0 0 0 gpi[27]
port 21 nsew signal input
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 gpi[28]
port 22 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 gpi[29]
port 23 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 gpi[2]
port 24 nsew signal input
flabel metal3 s 0 39448 800 39568 0 FreeSans 480 0 0 0 gpi[30]
port 25 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 gpi[31]
port 26 nsew signal input
flabel metal2 s 24490 40762 24546 41562 0 FreeSans 224 90 0 0 gpi[32]
port 27 nsew signal input
flabel metal2 s 6458 40762 6514 41562 0 FreeSans 224 90 0 0 gpi[33]
port 28 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 gpi[3]
port 29 nsew signal input
flabel metal2 s 15474 40762 15530 41562 0 FreeSans 224 90 0 0 gpi[4]
port 30 nsew signal input
flabel metal2 s 37370 40762 37426 41562 0 FreeSans 224 90 0 0 gpi[5]
port 31 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 gpi[6]
port 32 nsew signal input
flabel metal2 s 19982 40762 20038 41562 0 FreeSans 224 90 0 0 gpi[7]
port 33 nsew signal input
flabel metal2 s 39302 40762 39358 41562 0 FreeSans 224 90 0 0 gpi[8]
port 34 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gpi[9]
port 35 nsew signal input
flabel metal2 s 17406 40762 17462 41562 0 FreeSans 224 90 0 0 gpo[0]
port 36 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 gpo[10]
port 37 nsew signal tristate
flabel metal3 s 38618 10888 39418 11008 0 FreeSans 480 0 0 0 gpo[11]
port 38 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 gpo[12]
port 39 nsew signal tristate
flabel metal3 s 38618 15648 39418 15768 0 FreeSans 480 0 0 0 gpo[13]
port 40 nsew signal tristate
flabel metal2 s 18 40762 74 41562 0 FreeSans 224 90 0 0 gpo[14]
port 41 nsew signal tristate
flabel metal2 s 26422 40762 26478 41562 0 FreeSans 224 90 0 0 gpo[15]
port 42 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gpo[16]
port 43 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 gpo[17]
port 44 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 gpo[18]
port 45 nsew signal tristate
flabel metal2 s 21914 40762 21970 41562 0 FreeSans 224 90 0 0 gpo[19]
port 46 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 gpo[1]
port 47 nsew signal tristate
flabel metal3 s 38618 38768 39418 38888 0 FreeSans 480 0 0 0 gpo[20]
port 48 nsew signal tristate
flabel metal2 s 12898 40762 12954 41562 0 FreeSans 224 90 0 0 gpo[21]
port 49 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 gpo[22]
port 50 nsew signal tristate
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 gpo[23]
port 51 nsew signal tristate
flabel metal3 s 38618 36728 39418 36848 0 FreeSans 480 0 0 0 gpo[24]
port 52 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 gpo[25]
port 53 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 gpo[26]
port 54 nsew signal tristate
flabel metal3 s 38618 34008 39418 34128 0 FreeSans 480 0 0 0 gpo[27]
port 55 nsew signal tristate
flabel metal3 s 38618 1368 39418 1488 0 FreeSans 480 0 0 0 gpo[28]
port 56 nsew signal tristate
flabel metal2 s 9034 40762 9090 41562 0 FreeSans 224 90 0 0 gpo[29]
port 57 nsew signal tristate
flabel metal3 s 38618 20408 39418 20528 0 FreeSans 480 0 0 0 gpo[2]
port 58 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 gpo[30]
port 59 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 gpo[31]
port 60 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 gpo[32]
port 61 nsew signal tristate
flabel metal3 s 38618 22448 39418 22568 0 FreeSans 480 0 0 0 gpo[33]
port 62 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 gpo[3]
port 63 nsew signal tristate
flabel metal2 s 35438 40762 35494 41562 0 FreeSans 224 90 0 0 gpo[4]
port 64 nsew signal tristate
flabel metal2 s 32862 40762 32918 41562 0 FreeSans 224 90 0 0 gpo[5]
port 65 nsew signal tristate
flabel metal2 s 4526 40762 4582 41562 0 FreeSans 224 90 0 0 gpo[6]
port 66 nsew signal tristate
flabel metal2 s 10966 40762 11022 41562 0 FreeSans 224 90 0 0 gpo[7]
port 67 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 gpo[8]
port 68 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 gpo[9]
port 69 nsew signal tristate
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 nrst
port 70 nsew signal input
flabel metal3 s 38618 17688 39418 17808 0 FreeSans 480 0 0 0 store_en
port 71 nsew signal tristate
flabel metal4 s 4208 2128 4528 39216 0 FreeSans 1920 90 0 0 vccd1
port 72 nsew power bidirectional
flabel metal4 s 34928 2128 35248 39216 0 FreeSans 1920 90 0 0 vccd1
port 72 nsew power bidirectional
flabel metal4 s 19568 2128 19888 39216 0 FreeSans 1920 90 0 0 vssd1
port 73 nsew ground bidirectional
rlabel metal1 19688 38624 19688 38624 0 vccd1
rlabel via1 19688 39168 19688 39168 0 vssd1
rlabel metal1 19826 23732 19826 23732 0 ALU.flags_to_alu\[0\]
rlabel metal1 9522 33932 9522 33932 0 ALU.flags_to_alu\[1\]
rlabel metal2 8418 26622 8418 26622 0 ALU.flags_to_alu\[2\]
rlabel metal1 15410 29648 15410 29648 0 ALU.flags_to_alu\[3\]
rlabel metal1 18768 28118 18768 28118 0 ALU.flags_to_alu\[4\]
rlabel metal1 6670 31892 6670 31892 0 ALU.flags_to_alu\[5\]
rlabel metal1 10810 23834 10810 23834 0 ALU.flags_to_alu\[6\]
rlabel metal1 16100 34510 16100 34510 0 ALU.flags_to_alu\[7\]
rlabel metal2 9614 12920 9614 12920 0 ALU.immediate\[0\]
rlabel metal1 6348 13362 6348 13362 0 ALU.immediate\[10\]
rlabel metal2 16606 21488 16606 21488 0 ALU.immediate\[11\]
rlabel metal1 9246 18054 9246 18054 0 ALU.immediate\[12\]
rlabel metal1 7820 17850 7820 17850 0 ALU.immediate\[13\]
rlabel metal1 8096 12954 8096 12954 0 ALU.immediate\[14\]
rlabel metal2 17250 19924 17250 19924 0 ALU.immediate\[15\]
rlabel metal1 17802 7888 17802 7888 0 ALU.immediate\[1\]
rlabel metal1 17894 9146 17894 9146 0 ALU.immediate\[2\]
rlabel metal1 16836 8602 16836 8602 0 ALU.immediate\[3\]
rlabel metal2 21344 13940 21344 13940 0 ALU.immediate\[4\]
rlabel metal2 17618 11458 17618 11458 0 ALU.immediate\[5\]
rlabel metal1 11592 9146 11592 9146 0 ALU.immediate\[6\]
rlabel metal2 12282 16031 12282 16031 0 ALU.immediate\[7\]
rlabel metal1 13938 17136 13938 17136 0 ALU.immediate\[8\]
rlabel metal1 4462 19958 4462 19958 0 ALU.immediate\[9\]
rlabel metal1 13110 7174 13110 7174 0 ByteBuffer.counter\[0\]
rlabel metal1 13202 6834 13202 6834 0 ByteBuffer.counter\[1\]
rlabel metal1 12926 12818 12926 12818 0 ByteBuffer.instr\[16\]
rlabel metal1 15226 19788 15226 19788 0 ByteBuffer.instr\[17\]
rlabel metal2 16882 12614 16882 12614 0 ByteBuffer.instr\[18\]
rlabel metal1 13432 19754 13432 19754 0 ByteBuffer.instr\[19\]
rlabel metal1 15410 19822 15410 19822 0 ByteBuffer.instr\[20\]
rlabel metal1 19872 19754 19872 19754 0 ByteBuffer.instr\[21\]
rlabel metal1 13294 9588 13294 9588 0 ByteBuffer.instr\[22\]
rlabel metal2 15226 13090 15226 13090 0 ByteBuffer.instr\[23\]
rlabel metal1 11914 8466 11914 8466 0 ByteBuffer.next_counter\[0\]
rlabel metal2 9706 7514 9706 7514 0 ByteBuffer.next_counter\[1\]
rlabel metal2 8234 5372 8234 5372 0 ByteDecoder.num_bytes\[1\]
rlabel metal1 9982 5134 9982 5134 0 ByteDecoder.num_bytes\[2\]
rlabel metal1 9062 5780 9062 5780 0 ByteDecoder.num_bytes\[3\]
rlabel metal1 12696 5678 12696 5678 0 ByteDecoder.state\[0\]
rlabel metal1 12512 5678 12512 5678 0 ByteDecoder.state\[1\]
rlabel metal1 10304 5202 10304 5202 0 FSM.next_state\[0\]
rlabel metal1 11776 5270 11776 5270 0 FSM.next_state\[1\]
rlabel metal2 15410 6800 15410 6800 0 MemControl.state\[0\]
rlabel metal2 15870 4964 15870 4964 0 MemControl.state\[1\]
rlabel metal1 14858 6154 14858 6154 0 MemControl.state\[2\]
rlabel metal1 9614 8058 9614 8058 0 PC.i_mem_addr\[0\]
rlabel metal1 2530 23018 2530 23018 0 PC.i_mem_addr\[10\]
rlabel metal1 3910 20876 3910 20876 0 PC.i_mem_addr\[11\]
rlabel metal2 7958 22848 7958 22848 0 PC.i_mem_addr\[12\]
rlabel metal1 4922 24922 4922 24922 0 PC.i_mem_addr\[13\]
rlabel metal1 4416 24174 4416 24174 0 PC.i_mem_addr\[14\]
rlabel metal1 5152 19822 5152 19822 0 PC.i_mem_addr\[15\]
rlabel metal1 5796 7378 5796 7378 0 PC.i_mem_addr\[1\]
rlabel metal1 4462 8466 4462 8466 0 PC.i_mem_addr\[2\]
rlabel metal1 6624 10778 6624 10778 0 PC.i_mem_addr\[3\]
rlabel metal1 4324 12138 4324 12138 0 PC.i_mem_addr\[4\]
rlabel metal1 3588 12954 3588 12954 0 PC.i_mem_addr\[5\]
rlabel metal1 3358 14994 3358 14994 0 PC.i_mem_addr\[6\]
rlabel metal1 5842 17238 5842 17238 0 PC.i_mem_addr\[7\]
rlabel metal1 17388 14042 17388 14042 0 PC.i_mem_addr\[8\]
rlabel metal1 3680 20366 3680 20366 0 PC.i_mem_addr\[9\]
rlabel metal1 30406 25330 30406 25330 0 RegFile.A\[0\]
rlabel metal1 21942 33456 21942 33456 0 RegFile.A\[1\]
rlabel via2 18998 26979 18998 26979 0 RegFile.A\[2\]
rlabel metal1 18860 29138 18860 29138 0 RegFile.A\[3\]
rlabel metal2 13754 24327 13754 24327 0 RegFile.A\[4\]
rlabel metal2 32522 30464 32522 30464 0 RegFile.A\[5\]
rlabel metal2 13156 35564 13156 35564 0 RegFile.A\[6\]
rlabel metal1 36524 33898 36524 33898 0 RegFile.A\[7\]
rlabel metal1 28428 25194 28428 25194 0 RegFile.B\[0\]
rlabel metal1 20102 33898 20102 33898 0 RegFile.B\[1\]
rlabel metal1 15042 26452 15042 26452 0 RegFile.B\[2\]
rlabel metal1 17250 29512 17250 29512 0 RegFile.B\[3\]
rlabel metal2 30038 28832 30038 28832 0 RegFile.B\[4\]
rlabel viali 29670 31790 29670 31790 0 RegFile.B\[5\]
rlabel metal1 27186 37230 27186 37230 0 RegFile.B\[6\]
rlabel metal1 24150 35734 24150 35734 0 RegFile.B\[7\]
rlabel metal1 20746 25806 20746 25806 0 RegFile.C\[0\]
rlabel viali 12097 34578 12097 34578 0 RegFile.C\[1\]
rlabel metal1 16652 28458 16652 28458 0 RegFile.C\[2\]
rlabel metal2 16238 31246 16238 31246 0 RegFile.C\[3\]
rlabel metal1 19182 29784 19182 29784 0 RegFile.C\[4\]
rlabel metal2 20746 30957 20746 30957 0 RegFile.C\[5\]
rlabel metal1 11316 36142 11316 36142 0 RegFile.C\[6\]
rlabel metal2 21022 34884 21022 34884 0 RegFile.C\[7\]
rlabel metal1 22494 26928 22494 26928 0 RegFile.D\[0\]
rlabel metal2 33350 34816 33350 34816 0 RegFile.D\[1\]
rlabel metal1 16146 28560 16146 28560 0 RegFile.D\[2\]
rlabel metal2 16054 29308 16054 29308 0 RegFile.D\[3\]
rlabel via1 22016 29138 22016 29138 0 RegFile.D\[4\]
rlabel metal2 22034 31892 22034 31892 0 RegFile.D\[5\]
rlabel metal1 16008 37842 16008 37842 0 RegFile.D\[6\]
rlabel metal2 30038 35972 30038 35972 0 RegFile.D\[7\]
rlabel via1 13110 25466 13110 25466 0 RegFile.E\[0\]
rlabel metal1 7728 35802 7728 35802 0 RegFile.E\[1\]
rlabel metal1 14766 26248 14766 26248 0 RegFile.E\[2\]
rlabel metal1 14674 30668 14674 30668 0 RegFile.E\[3\]
rlabel metal1 16146 27608 16146 27608 0 RegFile.E\[4\]
rlabel metal2 6762 33728 6762 33728 0 RegFile.E\[5\]
rlabel metal2 16882 36992 16882 36992 0 RegFile.E\[6\]
rlabel metal1 24242 37774 24242 37774 0 RegFile.E\[7\]
rlabel metal1 22586 25160 22586 25160 0 RegFile.H\[0\]
rlabel metal1 26450 33966 26450 33966 0 RegFile.H\[1\]
rlabel metal1 25162 26282 25162 26282 0 RegFile.H\[2\]
rlabel metal2 17710 30515 17710 30515 0 RegFile.H\[3\]
rlabel metal1 26174 28526 26174 28526 0 RegFile.H\[4\]
rlabel metal2 32154 32572 32154 32572 0 RegFile.H\[5\]
rlabel metal2 25162 36176 25162 36176 0 RegFile.H\[6\]
rlabel metal1 33580 36142 33580 36142 0 RegFile.H\[7\]
rlabel metal1 12466 24752 12466 24752 0 RegFile.L\[0\]
rlabel metal1 8418 34476 8418 34476 0 RegFile.L\[1\]
rlabel via1 16790 28050 16790 28050 0 RegFile.L\[2\]
rlabel metal1 9430 30838 9430 30838 0 RegFile.L\[3\]
rlabel metal1 6026 29614 6026 29614 0 RegFile.L\[4\]
rlabel metal1 6440 32946 6440 32946 0 RegFile.L\[5\]
rlabel metal1 10672 37094 10672 37094 0 RegFile.L\[6\]
rlabel metal1 22540 37162 22540 37162 0 RegFile.L\[7\]
rlabel metal1 16652 4794 16652 4794 0 _0000_
rlabel metal1 13708 5270 13708 5270 0 _0001_
rlabel metal1 14536 4250 14536 4250 0 _0066_
rlabel metal1 7728 5746 7728 5746 0 _0067_
rlabel metal1 8326 4216 8326 4216 0 _0068_
rlabel metal1 6072 5338 6072 5338 0 _0069_
rlabel metal1 6578 15130 6578 15130 0 _0070_
rlabel metal1 6164 14042 6164 14042 0 _0071_
rlabel metal1 4830 12954 4830 12954 0 _0072_
rlabel metal1 6900 21114 6900 21114 0 _0073_
rlabel metal1 8004 17850 8004 17850 0 _0074_
rlabel metal1 6486 17306 6486 17306 0 _0075_
rlabel metal1 6440 12750 6440 12750 0 _0076_
rlabel metal1 6992 19482 6992 19482 0 _0077_
rlabel metal1 11270 13192 11270 13192 0 _0078_
rlabel metal1 13202 15130 13202 15130 0 _0079_
rlabel metal1 15170 12410 15170 12410 0 _0080_
rlabel metal1 11822 11696 11822 11696 0 _0081_
rlabel metal1 10212 14450 10212 14450 0 _0082_
rlabel metal1 14168 10710 14168 10710 0 _0083_
rlabel metal1 11822 9962 11822 9962 0 _0084_
rlabel metal1 13570 12886 13570 12886 0 _0085_
rlabel metal2 8602 13022 8602 13022 0 _0086_
rlabel metal1 15676 6970 15676 6970 0 _0087_
rlabel metal2 16054 9112 16054 9112 0 _0088_
rlabel metal1 13570 8398 13570 8398 0 _0089_
rlabel metal1 10258 11186 10258 11186 0 _0090_
rlabel metal1 16054 11186 16054 11186 0 _0091_
rlabel metal2 10074 9180 10074 9180 0 _0092_
rlabel metal1 9476 16218 9476 16218 0 _0093_
rlabel metal2 11086 22882 11086 22882 0 _0094_
rlabel metal1 7498 33082 7498 33082 0 _0095_
rlabel metal1 7360 26554 7360 26554 0 _0096_
rlabel metal1 5290 30158 5290 30158 0 _0097_
rlabel metal1 6532 28594 6532 28594 0 _0098_
rlabel metal1 5927 31994 5927 31994 0 _0099_
rlabel metal2 9338 23460 9338 23460 0 _0100_
rlabel metal1 5290 26010 5290 26010 0 _0101_
rlabel metal2 7958 24548 7958 24548 0 _0102_
rlabel metal1 7452 34714 7452 34714 0 _0103_
rlabel metal2 8326 27812 8326 27812 0 _0104_
rlabel metal2 8326 31552 8326 31552 0 _0105_
rlabel metal1 4600 28730 4600 28730 0 _0106_
rlabel metal1 4968 32538 4968 32538 0 _0107_
rlabel metal1 9246 37128 9246 37128 0 _0108_
rlabel metal1 20838 36890 20838 36890 0 _0109_
rlabel metal1 25944 24242 25944 24242 0 _0110_
rlabel metal1 31004 35122 31004 35122 0 _0111_
rlabel metal1 31372 26418 31372 26418 0 _0112_
rlabel metal2 35282 31450 35282 31450 0 _0113_
rlabel metal2 34454 28322 34454 28322 0 _0114_
rlabel metal1 31510 32776 31510 32776 0 _0115_
rlabel metal2 28198 35428 28198 35428 0 _0116_
rlabel metal2 32246 36516 32246 36516 0 _0117_
rlabel metal1 9016 25466 9016 25466 0 _0118_
rlabel metal1 6440 35802 6440 35802 0 _0119_
rlabel metal1 10166 27098 10166 27098 0 _0120_
rlabel metal1 6348 30362 6348 30362 0 _0121_
rlabel metal2 4646 27880 4646 27880 0 _0122_
rlabel metal1 5336 33898 5336 33898 0 _0123_
rlabel metal2 12834 38488 12834 38488 0 _0124_
rlabel metal1 21758 38216 21758 38216 0 _0125_
rlabel metal1 26542 27098 26542 27098 0 _0126_
rlabel metal1 33166 35122 33166 35122 0 _0127_
rlabel metal1 33534 26894 33534 26894 0 _0128_
rlabel metal1 34132 30906 34132 30906 0 _0129_
rlabel metal1 32246 28594 32246 28594 0 _0130_
rlabel metal1 28566 32538 28566 32538 0 _0131_
rlabel metal1 25944 37978 25944 37978 0 _0132_
rlabel metal1 30590 37298 30590 37298 0 _0133_
rlabel metal1 10580 24922 10580 24922 0 _0134_
rlabel metal1 9568 35734 9568 35734 0 _0135_
rlabel metal1 10580 28186 10580 28186 0 _0136_
rlabel metal1 9844 31450 9844 31450 0 _0137_
rlabel metal1 8878 29682 8878 29682 0 _0138_
rlabel metal1 9246 33592 9246 33592 0 _0139_
rlabel metal1 9706 37978 9706 37978 0 _0140_
rlabel metal1 19596 38386 19596 38386 0 _0141_
rlabel metal1 27876 26894 27876 26894 0 _0142_
rlabel metal2 28106 34272 28106 34272 0 _0143_
rlabel metal1 29762 27064 29762 27064 0 _0144_
rlabel metal1 27738 29206 27738 29206 0 _0145_
rlabel metal2 29302 28832 29302 28832 0 _0146_
rlabel metal1 28060 31654 28060 31654 0 _0147_
rlabel metal1 27186 37978 27186 37978 0 _0148_
rlabel metal1 29210 37774 29210 37774 0 _0149_
rlabel metal1 29026 24718 29026 24718 0 _0150_
rlabel metal1 34914 32946 34914 32946 0 _0151_
rlabel metal1 35098 26418 35098 26418 0 _0152_
rlabel metal1 34914 29002 34914 29002 0 _0153_
rlabel metal1 34776 25194 34776 25194 0 _0154_
rlabel metal1 30038 31246 30038 31246 0 _0155_
rlabel metal1 27048 33422 27048 33422 0 _0156_
rlabel metal1 34546 34034 34546 34034 0 _0157_
rlabel metal1 7452 7514 7452 7514 0 _0158_
rlabel metal1 4646 6426 4646 6426 0 _0159_
rlabel metal1 2944 7446 2944 7446 0 _0160_
rlabel metal1 4692 10234 4692 10234 0 _0161_
rlabel metal1 1748 10778 1748 10778 0 _0162_
rlabel metal1 1840 12410 1840 12410 0 _0163_
rlabel metal1 1840 14042 1840 14042 0 _0164_
rlabel metal2 4278 17442 4278 17442 0 _0165_
rlabel metal1 2024 16422 2024 16422 0 _0166_
rlabel metal1 1748 19414 1748 19414 0 _0167_
rlabel metal1 1748 24378 1748 24378 0 _0168_
rlabel metal1 1748 21590 1748 21590 0 _0169_
rlabel metal1 5612 24242 5612 24242 0 _0170_
rlabel metal1 3772 25466 3772 25466 0 _0171_
rlabel metal2 2898 25500 2898 25500 0 _0172_
rlabel metal1 4784 18938 4784 18938 0 _0173_
rlabel metal1 27968 4250 27968 4250 0 _0174_
rlabel metal1 27968 6698 27968 6698 0 _0175_
rlabel metal1 26082 8976 26082 8976 0 _0176_
rlabel metal1 26772 8466 26772 8466 0 _0177_
rlabel metal1 27554 6834 27554 6834 0 _0178_
rlabel viali 27554 6763 27554 6763 0 _0179_
rlabel metal1 28382 6732 28382 6732 0 _0180_
rlabel metal1 27922 7344 27922 7344 0 _0181_
rlabel metal1 28520 7378 28520 7378 0 _0182_
rlabel metal1 17664 10642 17664 10642 0 _0183_
rlabel metal1 36202 21658 36202 21658 0 _0184_
rlabel metal1 35650 20944 35650 20944 0 _0185_
rlabel metal1 35190 20876 35190 20876 0 _0186_
rlabel metal2 33350 20672 33350 20672 0 _0187_
rlabel metal2 33350 30328 33350 30328 0 _0188_
rlabel metal1 34592 29138 34592 29138 0 _0189_
rlabel metal2 23046 5644 23046 5644 0 _0190_
rlabel metal1 23368 5338 23368 5338 0 _0191_
rlabel metal1 23414 5100 23414 5100 0 _0192_
rlabel metal2 24426 4896 24426 4896 0 _0193_
rlabel metal1 20654 4794 20654 4794 0 _0194_
rlabel metal1 24886 5644 24886 5644 0 _0195_
rlabel metal1 25392 6426 25392 6426 0 _0196_
rlabel metal1 18952 8602 18952 8602 0 _0197_
rlabel metal1 25116 8806 25116 8806 0 _0198_
rlabel metal1 25392 7310 25392 7310 0 _0199_
rlabel metal1 25484 7446 25484 7446 0 _0200_
rlabel metal1 24610 5712 24610 5712 0 _0201_
rlabel metal1 24058 5134 24058 5134 0 _0202_
rlabel metal2 23690 5508 23690 5508 0 _0203_
rlabel metal1 14122 19244 14122 19244 0 _0204_
rlabel metal2 35926 19584 35926 19584 0 _0205_
rlabel metal1 35558 19890 35558 19890 0 _0206_
rlabel metal1 35374 19788 35374 19788 0 _0207_
rlabel metal1 34822 20026 34822 20026 0 _0208_
rlabel via1 25346 21590 25346 21590 0 _0209_
rlabel metal1 29578 26282 29578 26282 0 _0210_
rlabel metal1 34776 26010 34776 26010 0 _0211_
rlabel metal2 22034 7854 22034 7854 0 _0212_
rlabel metal1 22356 8262 22356 8262 0 _0213_
rlabel metal1 19964 6426 19964 6426 0 _0214_
rlabel metal1 20884 6834 20884 6834 0 _0215_
rlabel metal2 22402 7650 22402 7650 0 _0216_
rlabel metal1 20102 7820 20102 7820 0 _0217_
rlabel metal1 23552 8466 23552 8466 0 _0218_
rlabel metal1 22908 8942 22908 8942 0 _0219_
rlabel metal1 23230 8500 23230 8500 0 _0220_
rlabel metal1 22402 7854 22402 7854 0 _0221_
rlabel metal1 22448 7378 22448 7378 0 _0222_
rlabel metal1 23184 7514 23184 7514 0 _0223_
rlabel metal2 9062 19873 9062 19873 0 _0224_
rlabel metal1 34362 18190 34362 18190 0 _0225_
rlabel metal1 35190 18190 35190 18190 0 _0226_
rlabel metal1 34822 18326 34822 18326 0 _0227_
rlabel metal1 34040 17646 34040 17646 0 _0228_
rlabel metal2 17250 19040 17250 19040 0 _0229_
rlabel metal1 33718 34510 33718 34510 0 _0230_
rlabel metal1 34684 33490 34684 33490 0 _0231_
rlabel metal1 22126 10676 22126 10676 0 _0232_
rlabel metal1 21022 10166 21022 10166 0 _0233_
rlabel metal1 21022 10098 21022 10098 0 _0234_
rlabel metal1 21390 10132 21390 10132 0 _0235_
rlabel metal1 21390 10234 21390 10234 0 _0236_
rlabel metal1 22586 10098 22586 10098 0 _0237_
rlabel metal1 22448 9690 22448 9690 0 _0238_
rlabel metal1 21896 11118 21896 11118 0 _0239_
rlabel metal1 21758 11016 21758 11016 0 _0240_
rlabel metal2 22310 10642 22310 10642 0 _0241_
rlabel metal1 22586 10234 22586 10234 0 _0242_
rlabel metal2 10166 20145 10166 20145 0 _0243_
rlabel metal2 31878 17068 31878 17068 0 _0244_
rlabel metal1 32384 16762 32384 16762 0 _0245_
rlabel metal1 31878 17034 31878 17034 0 _0246_
rlabel metal1 33074 17136 33074 17136 0 _0247_
rlabel metal1 18676 14042 18676 14042 0 _0248_
rlabel metal1 26910 24854 26910 24854 0 _0249_
rlabel metal1 28980 23834 28980 23834 0 _0250_
rlabel metal1 24150 21658 24150 21658 0 _0251_
rlabel metal2 28382 24582 28382 24582 0 _0252_
rlabel metal1 29118 36890 29118 36890 0 _0253_
rlabel metal1 27002 37434 27002 37434 0 _0254_
rlabel metal1 28198 30906 28198 30906 0 _0255_
rlabel metal1 29348 28526 29348 28526 0 _0256_
rlabel metal1 28382 29614 28382 29614 0 _0257_
rlabel metal1 30176 26554 30176 26554 0 _0258_
rlabel metal1 28198 33966 28198 33966 0 _0259_
rlabel metal1 28014 26554 28014 26554 0 _0260_
rlabel metal1 13386 17510 13386 17510 0 _0261_
rlabel metal1 13570 21556 13570 21556 0 _0262_
rlabel metal1 13938 20026 13938 20026 0 _0263_
rlabel metal1 14720 21114 14720 21114 0 _0264_
rlabel metal1 23736 23698 23736 23698 0 _0265_
rlabel metal1 22586 21658 22586 21658 0 _0266_
rlabel metal2 22954 22916 22954 22916 0 _0267_
rlabel metal1 22724 23562 22724 23562 0 _0268_
rlabel metal1 22862 21930 22862 21930 0 _0269_
rlabel metal1 9614 33014 9614 33014 0 _0270_
rlabel metal2 19458 38454 19458 38454 0 _0271_
rlabel metal1 11270 37910 11270 37910 0 _0272_
rlabel metal1 10120 37842 10120 37842 0 _0273_
rlabel metal1 6302 32878 6302 32878 0 _0274_
rlabel metal1 10028 33082 10028 33082 0 _0275_
rlabel metal1 9568 21658 9568 21658 0 _0276_
rlabel metal1 8556 29274 8556 29274 0 _0277_
rlabel metal1 10028 20026 10028 20026 0 _0278_
rlabel metal1 10120 31314 10120 31314 0 _0279_
rlabel metal1 9660 21114 9660 21114 0 _0280_
rlabel metal1 11178 28050 11178 28050 0 _0281_
rlabel metal1 8280 34578 8280 34578 0 _0282_
rlabel metal1 9660 35258 9660 35258 0 _0283_
rlabel metal1 11132 19958 11132 19958 0 _0284_
rlabel metal1 11408 24786 11408 24786 0 _0285_
rlabel metal1 24978 23290 24978 23290 0 _0286_
rlabel metal2 25346 23970 25346 23970 0 _0287_
rlabel metal2 23506 24004 23506 24004 0 _0288_
rlabel via1 33166 27982 33166 27982 0 _0289_
rlabel metal1 31280 36890 31280 36890 0 _0290_
rlabel metal1 26266 37434 26266 37434 0 _0291_
rlabel metal1 29072 32402 29072 32402 0 _0292_
rlabel metal1 33028 28186 33028 28186 0 _0293_
rlabel metal1 33856 30702 33856 30702 0 _0294_
rlabel metal1 33212 26554 33212 26554 0 _0295_
rlabel metal1 33626 34714 33626 34714 0 _0296_
rlabel metal1 27002 26962 27002 26962 0 _0297_
rlabel metal1 23414 25908 23414 25908 0 _0298_
rlabel metal1 21666 37978 21666 37978 0 _0299_
rlabel metal1 12190 37978 12190 37978 0 _0300_
rlabel metal1 5520 33626 5520 33626 0 _0301_
rlabel metal1 5612 27438 5612 27438 0 _0302_
rlabel metal1 6946 30226 6946 30226 0 _0303_
rlabel metal1 11040 26962 11040 26962 0 _0304_
rlabel metal1 6831 35666 6831 35666 0 _0305_
rlabel metal1 9292 25262 9292 25262 0 _0306_
rlabel metal2 23966 23324 23966 23324 0 _0307_
rlabel metal1 31786 34476 31786 34476 0 _0308_
rlabel metal1 32338 36142 32338 36142 0 _0309_
rlabel metal1 28244 35054 28244 35054 0 _0310_
rlabel metal1 31096 32266 31096 32266 0 _0311_
rlabel metal1 34408 28050 34408 28050 0 _0312_
rlabel metal2 35466 31348 35466 31348 0 _0313_
rlabel metal1 31924 26010 31924 26010 0 _0314_
rlabel metal1 31326 34714 31326 34714 0 _0315_
rlabel metal1 26588 24786 26588 24786 0 _0316_
rlabel metal2 9890 36283 9890 36283 0 _0317_
rlabel metal1 21597 36754 21597 36754 0 _0318_
rlabel metal1 8832 36890 8832 36890 0 _0319_
rlabel metal1 5750 32402 5750 32402 0 _0320_
rlabel metal1 5106 28526 5106 28526 0 _0321_
rlabel metal1 8740 30906 8740 30906 0 _0322_
rlabel metal1 8510 27506 8510 27506 0 _0323_
rlabel metal1 7912 34578 7912 34578 0 _0324_
rlabel metal1 8142 24208 8142 24208 0 _0325_
rlabel metal2 6026 18785 6026 18785 0 _0326_
rlabel metal1 17802 20264 17802 20264 0 _0327_
rlabel metal1 11408 21658 11408 21658 0 _0328_
rlabel metal1 18124 18870 18124 18870 0 _0329_
rlabel metal2 18078 18122 18078 18122 0 _0330_
rlabel metal2 17710 18190 17710 18190 0 _0331_
rlabel metal1 15640 17714 15640 17714 0 _0332_
rlabel metal1 15272 17850 15272 17850 0 _0333_
rlabel via2 24334 23579 24334 23579 0 _0334_
rlabel metal1 8740 26418 8740 26418 0 _0335_
rlabel metal1 6302 25874 6302 25874 0 _0336_
rlabel metal2 9476 27540 9476 27540 0 _0337_
rlabel metal1 24702 20366 24702 20366 0 _0338_
rlabel metal1 24058 20026 24058 20026 0 _0339_
rlabel metal2 23874 19686 23874 19686 0 _0340_
rlabel metal1 22770 19482 22770 19482 0 _0341_
rlabel metal1 23644 19754 23644 19754 0 _0342_
rlabel metal2 23506 19737 23506 19737 0 _0343_
rlabel metal1 10028 22202 10028 22202 0 _0344_
rlabel metal1 9706 22746 9706 22746 0 _0345_
rlabel metal1 35742 15436 35742 15436 0 _0346_
rlabel metal1 28566 15028 28566 15028 0 _0347_
rlabel metal1 30084 7514 30084 7514 0 _0348_
rlabel metal2 33074 7378 33074 7378 0 _0349_
rlabel metal1 23966 6358 23966 6358 0 _0350_
rlabel metal1 24613 6426 24613 6426 0 _0351_
rlabel metal1 24150 7412 24150 7412 0 _0352_
rlabel metal2 24886 7004 24886 7004 0 _0353_
rlabel metal2 33166 6630 33166 6630 0 _0354_
rlabel metal1 34040 6630 34040 6630 0 _0355_
rlabel metal2 33534 10438 33534 10438 0 _0356_
rlabel metal1 33810 10438 33810 10438 0 _0357_
rlabel metal1 28842 10540 28842 10540 0 _0358_
rlabel metal1 34546 10506 34546 10506 0 _0359_
rlabel metal1 35374 10778 35374 10778 0 _0360_
rlabel metal1 34914 16626 34914 16626 0 _0361_
rlabel metal2 34546 18700 34546 18700 0 _0362_
rlabel metal1 34270 16966 34270 16966 0 _0363_
rlabel metal1 34316 17170 34316 17170 0 _0364_
rlabel metal1 34914 16490 34914 16490 0 _0365_
rlabel metal1 35236 16762 35236 16762 0 _0366_
rlabel metal1 33994 15028 33994 15028 0 _0367_
rlabel metal1 31142 14382 31142 14382 0 _0368_
rlabel metal1 32476 14586 32476 14586 0 _0369_
rlabel metal1 33442 14892 33442 14892 0 _0370_
rlabel metal1 34592 15130 34592 15130 0 _0371_
rlabel metal1 35190 16048 35190 16048 0 _0372_
rlabel metal1 35236 15878 35236 15878 0 _0373_
rlabel metal1 34914 16694 34914 16694 0 _0374_
rlabel metal1 35098 16456 35098 16456 0 _0375_
rlabel metal1 29394 17034 29394 17034 0 _0376_
rlabel metal1 28704 17238 28704 17238 0 _0377_
rlabel metal1 28244 17034 28244 17034 0 _0378_
rlabel metal2 28382 17476 28382 17476 0 _0379_
rlabel metal1 22770 17170 22770 17170 0 _0380_
rlabel metal1 25254 17714 25254 17714 0 _0381_
rlabel metal1 25070 17714 25070 17714 0 _0382_
rlabel metal1 25944 17646 25944 17646 0 _0383_
rlabel metal1 26312 17714 26312 17714 0 _0384_
rlabel metal1 27002 17748 27002 17748 0 _0385_
rlabel metal1 27692 17850 27692 17850 0 _0386_
rlabel metal2 27922 17850 27922 17850 0 _0387_
rlabel metal3 17204 17884 17204 17884 0 _0388_
rlabel metal1 8970 21862 8970 21862 0 _0389_
rlabel metal1 7958 26282 7958 26282 0 _0390_
rlabel metal1 8280 32946 8280 32946 0 _0391_
rlabel metal1 30360 16218 30360 16218 0 _0392_
rlabel metal1 29670 16762 29670 16762 0 _0393_
rlabel metal1 29670 12614 29670 12614 0 _0394_
rlabel metal1 22954 12308 22954 12308 0 _0395_
rlabel metal1 26680 12138 26680 12138 0 _0396_
rlabel metal1 25802 11866 25802 11866 0 _0397_
rlabel metal1 29670 12410 29670 12410 0 _0398_
rlabel metal1 29026 17204 29026 17204 0 _0399_
rlabel metal1 28658 19788 28658 19788 0 _0400_
rlabel metal1 28934 19278 28934 19278 0 _0401_
rlabel metal1 29210 19380 29210 19380 0 _0402_
rlabel metal1 29624 17170 29624 17170 0 _0403_
rlabel metal1 16606 17000 16606 17000 0 _0404_
rlabel metal1 12098 22202 12098 22202 0 _0405_
rlabel metal1 11408 22610 11408 22610 0 _0406_
rlabel metal2 7222 13600 7222 13600 0 _0407_
rlabel metal2 12374 7378 12374 7378 0 _0408_
rlabel metal1 15502 9486 15502 9486 0 _0409_
rlabel metal1 14398 7310 14398 7310 0 _0410_
rlabel metal1 16054 13158 16054 13158 0 _0411_
rlabel metal1 14582 6324 14582 6324 0 _0412_
rlabel metal2 13616 21454 13616 21454 0 _0413_
rlabel metal1 9706 5576 9706 5576 0 _0414_
rlabel metal2 9430 6018 9430 6018 0 _0415_
rlabel metal1 9798 5202 9798 5202 0 _0416_
rlabel metal1 13064 19686 13064 19686 0 _0417_
rlabel metal2 13202 20026 13202 20026 0 _0418_
rlabel metal1 8280 9622 8280 9622 0 _0419_
rlabel metal1 8924 14790 8924 14790 0 _0420_
rlabel metal1 14674 11118 14674 11118 0 _0421_
rlabel metal1 11362 15062 11362 15062 0 _0422_
rlabel metal1 8602 10608 8602 10608 0 _0423_
rlabel metal1 9246 10778 9246 10778 0 _0424_
rlabel metal1 8096 9554 8096 9554 0 _0425_
rlabel metal2 9522 14042 9522 14042 0 _0426_
rlabel metal1 7682 11152 7682 11152 0 _0427_
rlabel metal1 7912 11118 7912 11118 0 _0428_
rlabel metal1 8464 13226 8464 13226 0 _0429_
rlabel metal1 7820 9554 7820 9554 0 _0430_
rlabel metal1 7728 6222 7728 6222 0 _0431_
rlabel metal1 8326 6290 8326 6290 0 _0432_
rlabel metal1 9568 10098 9568 10098 0 _0433_
rlabel metal1 7958 9894 7958 9894 0 _0434_
rlabel metal2 15456 12818 15456 12818 0 _0435_
rlabel metal1 13570 14246 13570 14246 0 _0436_
rlabel metal1 9062 10132 9062 10132 0 _0437_
rlabel metal1 9338 6766 9338 6766 0 _0438_
rlabel metal1 9200 5202 9200 5202 0 _0439_
rlabel metal1 14398 18802 14398 18802 0 _0440_
rlabel metal1 14490 18292 14490 18292 0 _0441_
rlabel metal1 19550 18360 19550 18360 0 _0442_
rlabel metal1 16468 4590 16468 4590 0 _0443_
rlabel metal1 16100 4522 16100 4522 0 _0444_
rlabel metal1 2162 18156 2162 18156 0 _0445_
rlabel metal2 15042 12716 15042 12716 0 _0446_
rlabel metal1 36386 32538 36386 32538 0 _0447_
rlabel metal1 37030 18258 37030 18258 0 _0448_
rlabel metal1 9706 32946 9706 32946 0 _0449_
rlabel via3 12581 4012 12581 4012 0 _0450_
rlabel metal3 13271 4012 13271 4012 0 _0451_
rlabel metal1 1978 23800 1978 23800 0 _0452_
rlabel metal1 37352 28050 37352 28050 0 _0453_
rlabel metal1 2162 17646 2162 17646 0 _0454_
rlabel metal1 10994 8602 10994 8602 0 _0455_
rlabel metal1 14306 8908 14306 8908 0 _0456_
rlabel metal1 6532 9146 6532 9146 0 _0457_
rlabel metal1 4370 8976 4370 8976 0 _0458_
rlabel metal1 12190 10608 12190 10608 0 _0459_
rlabel metal1 3450 9588 3450 9588 0 _0460_
rlabel metal1 6670 13498 6670 13498 0 _0461_
rlabel metal2 3450 17476 3450 17476 0 _0462_
rlabel metal1 16606 16728 16606 16728 0 _0463_
rlabel metal2 17434 11084 17434 11084 0 _0464_
rlabel metal1 17250 3094 17250 3094 0 _0465_
rlabel metal1 1886 17646 1886 17646 0 _0466_
rlabel metal2 1978 4963 1978 4963 0 _0467_
rlabel metal2 2714 22916 2714 22916 0 _0468_
rlabel via2 5658 20859 5658 20859 0 _0469_
rlabel metal1 24840 21998 24840 21998 0 _0470_
rlabel metal2 12558 22780 12558 22780 0 _0471_
rlabel metal1 5934 21488 5934 21488 0 _0472_
rlabel metal1 2346 18326 2346 18326 0 _0473_
rlabel metal2 2530 17307 2530 17307 0 _0474_
rlabel metal2 27738 21760 27738 21760 0 _0475_
rlabel metal1 25530 37774 25530 37774 0 _0476_
rlabel metal1 20562 38454 20562 38454 0 _0477_
rlabel metal2 2162 16286 2162 16286 0 _0478_
rlabel metal1 37214 20842 37214 20842 0 _0479_
rlabel metal1 23000 3026 23000 3026 0 _0480_
rlabel metal1 34730 38250 34730 38250 0 _0481_
rlabel metal1 29394 37638 29394 37638 0 _0482_
rlabel metal2 5198 38369 5198 38369 0 _0483_
rlabel via2 12558 37859 12558 37859 0 _0484_
rlabel metal2 14398 4828 14398 4828 0 _0485_
rlabel metal1 7038 5202 7038 5202 0 _0486_
rlabel metal1 6992 14994 6992 14994 0 _0487_
rlabel metal1 6624 13906 6624 13906 0 _0488_
rlabel metal1 5520 12818 5520 12818 0 _0489_
rlabel metal1 13110 11050 13110 11050 0 _0490_
rlabel metal1 7176 20910 7176 20910 0 _0491_
rlabel metal1 8602 17646 8602 17646 0 _0492_
rlabel metal1 6854 17170 6854 17170 0 _0493_
rlabel metal1 6026 12852 6026 12852 0 _0494_
rlabel metal1 7222 19414 7222 19414 0 _0495_
rlabel metal1 13294 8058 13294 8058 0 _0496_
rlabel metal1 12788 13362 12788 13362 0 _0497_
rlabel metal1 10948 13226 10948 13226 0 _0498_
rlabel metal1 13800 14586 13800 14586 0 _0499_
rlabel metal2 15088 12580 15088 12580 0 _0500_
rlabel metal2 12006 11526 12006 11526 0 _0501_
rlabel metal1 11040 14994 11040 14994 0 _0502_
rlabel metal1 13938 11118 13938 11118 0 _0503_
rlabel metal1 11638 9690 11638 9690 0 _0504_
rlabel metal1 13708 13294 13708 13294 0 _0505_
rlabel metal1 8970 13294 8970 13294 0 _0506_
rlabel metal1 15456 7378 15456 7378 0 _0507_
rlabel metal1 16100 9554 16100 9554 0 _0508_
rlabel metal1 13156 8466 13156 8466 0 _0509_
rlabel metal1 9798 11220 9798 11220 0 _0510_
rlabel metal2 15594 11322 15594 11322 0 _0511_
rlabel metal1 10304 9554 10304 9554 0 _0512_
rlabel metal1 9752 16082 9752 16082 0 _0513_
rlabel metal1 17848 26010 17848 26010 0 _0514_
rlabel metal2 19090 30753 19090 30753 0 _0515_
rlabel via2 21298 32419 21298 32419 0 _0516_
rlabel via2 21298 31773 21298 31773 0 _0517_
rlabel metal1 18354 16150 18354 16150 0 _0518_
rlabel metal1 17434 7854 17434 7854 0 _0519_
rlabel metal1 10488 13498 10488 13498 0 _0520_
rlabel metal1 10304 12818 10304 12818 0 _0521_
rlabel metal1 10120 8602 10120 8602 0 _0522_
rlabel metal1 11454 18258 11454 18258 0 _0523_
rlabel metal1 12696 17850 12696 17850 0 _0524_
rlabel metal2 12558 17459 12558 17459 0 _0525_
rlabel metal1 11822 17646 11822 17646 0 _0526_
rlabel metal1 12466 17272 12466 17272 0 _0527_
rlabel metal2 12006 17510 12006 17510 0 _0528_
rlabel metal1 11546 17850 11546 17850 0 _0529_
rlabel metal2 11914 19788 11914 19788 0 _0530_
rlabel metal1 12650 19312 12650 19312 0 _0531_
rlabel metal1 12006 19414 12006 19414 0 _0532_
rlabel metal1 12190 18326 12190 18326 0 _0533_
rlabel metal1 11040 17714 11040 17714 0 _0534_
rlabel metal1 11132 18666 11132 18666 0 _0535_
rlabel metal1 11132 18734 11132 18734 0 _0536_
rlabel metal1 10396 17646 10396 17646 0 _0537_
rlabel metal1 12650 17714 12650 17714 0 _0538_
rlabel metal1 10810 17170 10810 17170 0 _0539_
rlabel metal1 10304 17714 10304 17714 0 _0540_
rlabel metal1 9108 8602 9108 8602 0 _0541_
rlabel metal2 13202 9486 13202 9486 0 _0542_
rlabel metal1 7958 7378 7958 7378 0 _0543_
rlabel metal1 17618 7786 17618 7786 0 _0544_
rlabel metal1 6486 7956 6486 7956 0 _0545_
rlabel metal1 6486 7310 6486 7310 0 _0546_
rlabel metal1 5888 7514 5888 7514 0 _0547_
rlabel metal1 5060 6290 5060 6290 0 _0548_
rlabel metal1 5474 8398 5474 8398 0 _0549_
rlabel metal1 5888 7854 5888 7854 0 _0550_
rlabel metal1 6210 10064 6210 10064 0 _0551_
rlabel metal1 5612 8058 5612 8058 0 _0552_
rlabel metal1 4692 8602 4692 8602 0 _0553_
rlabel metal1 3634 8466 3634 8466 0 _0554_
rlabel metal2 13110 9962 13110 9962 0 _0555_
rlabel metal1 3713 12070 3713 12070 0 _0556_
rlabel metal2 6210 10438 6210 10438 0 _0557_
rlabel metal1 6486 10574 6486 10574 0 _0558_
rlabel metal1 5658 10132 5658 10132 0 _0559_
rlabel metal1 5014 10030 5014 10030 0 _0560_
rlabel metal1 10028 10438 10028 10438 0 _0561_
rlabel metal1 3726 10642 3726 10642 0 _0562_
rlabel metal1 3312 10778 3312 10778 0 _0563_
rlabel metal1 2162 10642 2162 10642 0 _0564_
rlabel metal1 18400 12138 18400 12138 0 _0565_
rlabel metal1 15042 12308 15042 12308 0 _0566_
rlabel metal1 4646 12750 4646 12750 0 _0567_
rlabel metal2 4554 12818 4554 12818 0 _0568_
rlabel metal1 4324 12886 4324 12886 0 _0569_
rlabel metal1 3358 12614 3358 12614 0 _0570_
rlabel metal1 2392 12206 2392 12206 0 _0571_
rlabel metal1 4784 15130 4784 15130 0 _0572_
rlabel metal1 4554 15572 4554 15572 0 _0573_
rlabel metal1 3864 14382 3864 14382 0 _0574_
rlabel metal2 4094 14722 4094 14722 0 _0575_
rlabel metal1 3358 15130 3358 15130 0 _0576_
rlabel metal1 2346 13906 2346 13906 0 _0577_
rlabel metal1 8740 15946 8740 15946 0 _0578_
rlabel metal1 5336 15674 5336 15674 0 _0579_
rlabel metal1 5106 16218 5106 16218 0 _0580_
rlabel metal1 4508 17170 4508 17170 0 _0581_
rlabel metal1 3588 19346 3588 19346 0 _0582_
rlabel metal1 4094 16456 4094 16456 0 _0583_
rlabel metal1 3910 15674 3910 15674 0 _0584_
rlabel metal1 9706 19856 9706 19856 0 _0585_
rlabel metal1 2806 16660 2806 16660 0 _0586_
rlabel metal1 2346 16490 2346 16490 0 _0587_
rlabel metal1 3964 21862 3964 21862 0 _0588_
rlabel metal1 4094 19788 4094 19788 0 _0589_
rlabel metal2 3910 19618 3910 19618 0 _0590_
rlabel metal1 3358 20026 3358 20026 0 _0591_
rlabel metal1 2208 19822 2208 19822 0 _0592_
rlabel metal2 4002 22848 4002 22848 0 _0593_
rlabel metal1 3312 22746 3312 22746 0 _0594_
rlabel metal1 2898 23290 2898 23290 0 _0595_
rlabel metal1 2162 24174 2162 24174 0 _0596_
rlabel metal1 4232 21998 4232 21998 0 _0597_
rlabel metal1 4370 21590 4370 21590 0 _0598_
rlabel metal1 4508 21114 4508 21114 0 _0599_
rlabel metal1 3910 21522 3910 21522 0 _0600_
rlabel metal2 1978 21828 1978 21828 0 _0601_
rlabel metal1 7314 22984 7314 22984 0 _0602_
rlabel viali 7223 23058 7223 23058 0 _0603_
rlabel metal2 7038 23494 7038 23494 0 _0604_
rlabel metal1 6164 23834 6164 23834 0 _0605_
rlabel metal1 5980 23290 5980 23290 0 _0606_
rlabel metal2 5290 23256 5290 23256 0 _0607_
rlabel metal1 5198 23120 5198 23120 0 _0608_
rlabel metal1 4922 23290 4922 23290 0 _0609_
rlabel metal2 4370 25092 4370 25092 0 _0610_
rlabel metal1 5382 22746 5382 22746 0 _0611_
rlabel metal1 4784 22746 4784 22746 0 _0612_
rlabel metal1 4462 23290 4462 23290 0 _0613_
rlabel metal1 3450 24378 3450 24378 0 _0614_
rlabel metal1 6394 19890 6394 19890 0 _0615_
rlabel metal1 5842 19686 5842 19686 0 _0616_
rlabel metal1 5060 18734 5060 18734 0 _0617_
rlabel metal1 17894 17612 17894 17612 0 _0618_
rlabel metal2 20010 17442 20010 17442 0 _0619_
rlabel metal1 18538 18666 18538 18666 0 _0620_
rlabel metal1 16422 17680 16422 17680 0 _0621_
rlabel metal1 19826 21522 19826 21522 0 _0622_
rlabel metal1 14306 22644 14306 22644 0 _0623_
rlabel metal1 14536 17102 14536 17102 0 _0624_
rlabel metal1 15364 13498 15364 13498 0 _0625_
rlabel metal1 19412 21522 19412 21522 0 _0626_
rlabel metal1 14260 15674 14260 15674 0 _0627_
rlabel metal1 13754 17680 13754 17680 0 _0628_
rlabel metal2 20654 33439 20654 33439 0 _0629_
rlabel metal1 29026 19380 29026 19380 0 _0630_
rlabel metal1 23966 18870 23966 18870 0 _0631_
rlabel metal1 15501 21556 15501 21556 0 _0632_
rlabel metal1 15870 20570 15870 20570 0 _0633_
rlabel metal2 15502 21556 15502 21556 0 _0634_
rlabel metal1 15739 16490 15739 16490 0 _0635_
rlabel metal1 11960 19210 11960 19210 0 _0636_
rlabel metal1 15226 20570 15226 20570 0 _0637_
rlabel metal1 14444 22066 14444 22066 0 _0638_
rlabel metal2 15594 17680 15594 17680 0 _0639_
rlabel metal1 15129 21556 15129 21556 0 _0640_
rlabel metal1 19412 20230 19412 20230 0 _0641_
rlabel metal1 18906 20774 18906 20774 0 _0642_
rlabel metal1 16284 19346 16284 19346 0 _0643_
rlabel metal1 16606 21998 16606 21998 0 _0644_
rlabel metal2 13386 14178 13386 14178 0 _0645_
rlabel metal1 16514 21862 16514 21862 0 _0646_
rlabel metal1 16744 17646 16744 17646 0 _0647_
rlabel metal1 16514 17578 16514 17578 0 _0648_
rlabel metal1 20792 18938 20792 18938 0 _0649_
rlabel metal2 20470 22916 20470 22916 0 _0650_
rlabel metal2 20838 23494 20838 23494 0 _0651_
rlabel metal1 21252 23766 21252 23766 0 _0652_
rlabel metal1 14168 23290 14168 23290 0 _0653_
rlabel metal1 18446 27472 18446 27472 0 _0654_
rlabel metal1 18538 17646 18538 17646 0 _0655_
rlabel metal1 17066 14416 17066 14416 0 _0656_
rlabel metal2 17066 14790 17066 14790 0 _0657_
rlabel metal1 12512 6290 12512 6290 0 _0658_
rlabel metal1 12834 21862 12834 21862 0 _0659_
rlabel metal1 16376 15470 16376 15470 0 _0660_
rlabel metal2 16698 16864 16698 16864 0 _0661_
rlabel metal1 16652 14382 16652 14382 0 _0662_
rlabel metal1 16238 14586 16238 14586 0 _0663_
rlabel metal1 18216 14926 18216 14926 0 _0664_
rlabel metal1 19918 19890 19918 19890 0 _0665_
rlabel metal1 19090 15436 19090 15436 0 _0666_
rlabel metal1 19412 18394 19412 18394 0 _0667_
rlabel metal1 18722 18734 18722 18734 0 _0668_
rlabel metal1 18630 16082 18630 16082 0 _0669_
rlabel metal1 18906 21114 18906 21114 0 _0670_
rlabel metal2 18262 16524 18262 16524 0 _0671_
rlabel metal2 18170 16252 18170 16252 0 _0672_
rlabel metal1 18722 15538 18722 15538 0 _0673_
rlabel metal1 18584 11050 18584 11050 0 _0674_
rlabel metal1 18906 15640 18906 15640 0 _0675_
rlabel metal1 30360 28934 30360 28934 0 _0676_
rlabel metal1 14904 23698 14904 23698 0 _0677_
rlabel metal1 20378 14960 20378 14960 0 _0678_
rlabel metal1 13892 21590 13892 21590 0 _0679_
rlabel viali 27648 25262 27648 25262 0 _0680_
rlabel metal1 13432 33966 13432 33966 0 _0681_
rlabel metal1 13662 35734 13662 35734 0 _0682_
rlabel viali 12192 32878 12192 32878 0 _0683_
rlabel metal1 19918 23664 19918 23664 0 _0684_
rlabel metal1 11730 36006 11730 36006 0 _0685_
rlabel metal1 14674 24378 14674 24378 0 _0686_
rlabel metal1 12236 34578 12236 34578 0 _0687_
rlabel metal1 28106 36346 28106 36346 0 _0688_
rlabel metal3 29233 33116 29233 33116 0 _0689_
rlabel metal2 30222 23324 30222 23324 0 _0690_
rlabel metal1 30498 22576 30498 22576 0 _0691_
rlabel metal1 18814 15334 18814 15334 0 _0692_
rlabel metal1 18262 16660 18262 16660 0 _0693_
rlabel metal1 17342 22576 17342 22576 0 _0694_
rlabel metal2 18722 19924 18722 19924 0 _0695_
rlabel metal1 18170 19754 18170 19754 0 _0696_
rlabel metal1 13432 19890 13432 19890 0 _0697_
rlabel metal2 17158 22848 17158 22848 0 _0698_
rlabel metal1 16054 32878 16054 32878 0 _0699_
rlabel metal1 17618 21658 17618 21658 0 _0700_
rlabel metal2 20194 21828 20194 21828 0 _0701_
rlabel metal2 19458 20196 19458 20196 0 _0702_
rlabel metal1 16100 31790 16100 31790 0 _0703_
rlabel metal1 18722 31858 18722 31858 0 _0704_
rlabel metal1 17549 28050 17549 28050 0 _0705_
rlabel metal1 21666 32402 21666 32402 0 _0706_
rlabel metal1 16974 28016 16974 28016 0 _0707_
rlabel metal1 20746 33966 20746 33966 0 _0708_
rlabel metal2 17066 36380 17066 36380 0 _0709_
rlabel metal1 26266 35632 26266 35632 0 _0710_
rlabel metal2 20838 26180 20838 26180 0 _0711_
rlabel metal1 26542 35088 26542 35088 0 _0712_
rlabel metal1 26082 35156 26082 35156 0 _0713_
rlabel metal1 29670 22644 29670 22644 0 _0714_
rlabel metal1 30636 20434 30636 20434 0 _0715_
rlabel metal1 29624 22406 29624 22406 0 _0716_
rlabel metal1 30130 22746 30130 22746 0 _0717_
rlabel metal1 30222 22066 30222 22066 0 _0718_
rlabel metal1 31786 29172 31786 29172 0 _0719_
rlabel metal1 32062 29138 32062 29138 0 _0720_
rlabel metal1 34730 23188 34730 23188 0 _0721_
rlabel metal1 26726 29682 26726 29682 0 _0722_
rlabel metal1 25990 29648 25990 29648 0 _0723_
rlabel metal1 25668 29478 25668 29478 0 _0724_
rlabel metal1 27554 21080 27554 21080 0 _0725_
rlabel metal1 35282 21522 35282 21522 0 _0726_
rlabel metal2 31786 26588 31786 26588 0 _0727_
rlabel metal1 32982 25908 32982 25908 0 _0728_
rlabel metal1 35144 23086 35144 23086 0 _0729_
rlabel metal1 26542 26384 26542 26384 0 _0730_
rlabel metal1 26128 25874 26128 25874 0 _0731_
rlabel metal1 26956 22066 26956 22066 0 _0732_
rlabel metal2 27554 22984 27554 22984 0 _0733_
rlabel metal1 36754 22066 36754 22066 0 _0734_
rlabel metal1 36892 21998 36892 21998 0 _0735_
rlabel metal1 35880 22066 35880 22066 0 _0736_
rlabel metal1 36294 20026 36294 20026 0 _0737_
rlabel metal1 31786 34000 31786 34000 0 _0738_
rlabel metal1 32338 32402 32338 32402 0 _0739_
rlabel metal1 33212 19822 33212 19822 0 _0740_
rlabel metal1 20930 33354 20930 33354 0 _0741_
rlabel metal1 25898 34000 25898 34000 0 _0742_
rlabel metal1 25254 33320 25254 33320 0 _0743_
rlabel metal2 25346 20485 25346 20485 0 _0744_
rlabel metal1 33626 19856 33626 19856 0 _0745_
rlabel metal1 34868 19346 34868 19346 0 _0746_
rlabel metal1 28750 25296 28750 25296 0 _0747_
rlabel metal1 30038 25228 30038 25228 0 _0748_
rlabel metal1 31280 18734 31280 18734 0 _0749_
rlabel metal1 25254 25228 25254 25228 0 _0750_
rlabel metal2 24794 25670 24794 25670 0 _0751_
rlabel via3 25277 37332 25277 37332 0 _0752_
rlabel metal1 31004 18258 31004 18258 0 _0753_
rlabel metal1 31947 18326 31947 18326 0 _0754_
rlabel metal1 31464 18258 31464 18258 0 _0755_
rlabel metal1 32844 18326 32844 18326 0 _0756_
rlabel metal1 17204 19958 17204 19958 0 _0757_
rlabel metal1 17848 21522 17848 21522 0 _0758_
rlabel metal2 17434 22372 17434 22372 0 _0759_
rlabel metal1 13662 33830 13662 33830 0 _0760_
rlabel via2 14306 23749 14306 23749 0 _0761_
rlabel metal1 14168 33626 14168 33626 0 _0762_
rlabel metal2 15594 35207 15594 35207 0 _0763_
rlabel metal2 22862 31756 22862 31756 0 _0764_
rlabel metal1 15870 24242 15870 24242 0 _0765_
rlabel metal1 19734 24208 19734 24208 0 _0766_
rlabel metal1 14398 33932 14398 33932 0 _0767_
rlabel metal1 21620 30906 21620 30906 0 _0768_
rlabel metal1 22770 31246 22770 31246 0 _0769_
rlabel metal1 15778 36584 15778 36584 0 _0770_
rlabel metal2 17894 24922 17894 24922 0 _0771_
rlabel metal1 15732 23834 15732 23834 0 _0772_
rlabel via2 23046 31331 23046 31331 0 _0773_
rlabel metal1 20792 33490 20792 33490 0 _0774_
rlabel metal1 22908 18938 22908 18938 0 _0775_
rlabel metal2 12374 32640 12374 32640 0 _0776_
rlabel metal1 12190 32470 12190 32470 0 _0777_
rlabel metal3 14697 32028 14697 32028 0 _0778_
rlabel metal1 19044 11118 19044 11118 0 _0779_
rlabel metal1 18308 13226 18308 13226 0 _0780_
rlabel metal1 27324 8942 27324 8942 0 _0781_
rlabel via2 18722 11611 18722 11611 0 _0782_
rlabel metal1 18354 21114 18354 21114 0 _0783_
rlabel metal1 19506 36142 19506 36142 0 _0784_
rlabel metal1 17020 21114 17020 21114 0 _0785_
rlabel metal1 16284 28526 16284 28526 0 _0786_
rlabel metal1 25438 31824 25438 31824 0 _0787_
rlabel metal1 18492 37230 18492 37230 0 _0788_
rlabel metal2 20194 26792 20194 26792 0 _0789_
rlabel metal2 23966 32606 23966 32606 0 _0790_
rlabel metal2 25346 31994 25346 31994 0 _0791_
rlabel metal2 19090 31867 19090 31867 0 _0792_
rlabel metal2 20838 30141 20838 30141 0 _0793_
rlabel metal2 17710 33031 17710 33031 0 _0794_
rlabel metal1 22862 31450 22862 31450 0 _0795_
rlabel metal1 25162 31926 25162 31926 0 _0796_
rlabel metal1 25024 30906 25024 30906 0 _0797_
rlabel metal2 25622 31484 25622 31484 0 _0798_
rlabel metal1 20792 31314 20792 31314 0 _0799_
rlabel metal1 20976 31314 20976 31314 0 _0800_
rlabel metal1 22586 31144 22586 31144 0 _0801_
rlabel via3 26749 30396 26749 30396 0 _0802_
rlabel metal1 32338 10676 32338 10676 0 _0803_
rlabel metal1 32338 11152 32338 11152 0 _0804_
rlabel metal1 33442 13260 33442 13260 0 _0805_
rlabel metal2 33074 8704 33074 8704 0 _0806_
rlabel metal2 14674 27778 14674 27778 0 _0807_
rlabel metal1 14352 27914 14352 27914 0 _0808_
rlabel metal1 14260 26962 14260 26962 0 _0809_
rlabel metal2 15134 26656 15134 26656 0 _0810_
rlabel metal1 14582 26554 14582 26554 0 _0811_
rlabel metal1 14076 26554 14076 26554 0 _0812_
rlabel metal1 13570 26384 13570 26384 0 _0813_
rlabel metal2 13662 27098 13662 27098 0 _0814_
rlabel metal2 15824 21998 15824 21998 0 _0815_
rlabel metal1 18354 8908 18354 8908 0 _0816_
rlabel metal2 21114 34850 21114 34850 0 _0817_
rlabel metal2 16698 27268 16698 27268 0 _0818_
rlabel metal2 17802 27132 17802 27132 0 _0819_
rlabel metal1 16744 26282 16744 26282 0 _0820_
rlabel metal1 17572 26554 17572 26554 0 _0821_
rlabel metal1 16606 28390 16606 28390 0 _0822_
rlabel metal1 18308 27098 18308 27098 0 _0823_
rlabel metal1 18722 27098 18722 27098 0 _0824_
rlabel metal2 16054 27846 16054 27846 0 _0825_
rlabel metal2 17434 27302 17434 27302 0 _0826_
rlabel metal1 18354 27404 18354 27404 0 _0827_
rlabel metal1 17480 15674 17480 15674 0 _0828_
rlabel metal2 16422 12852 16422 12852 0 _0829_
rlabel metal2 18078 10234 18078 10234 0 _0830_
rlabel metal1 19918 4658 19918 4658 0 _0831_
rlabel metal1 30268 5202 30268 5202 0 _0832_
rlabel metal1 16652 29818 16652 29818 0 _0833_
rlabel metal1 17526 30158 17526 30158 0 _0834_
rlabel metal1 17066 30906 17066 30906 0 _0835_
rlabel metal2 17894 30566 17894 30566 0 _0836_
rlabel metal1 17112 30226 17112 30226 0 _0837_
rlabel metal1 18630 29648 18630 29648 0 _0838_
rlabel metal1 18814 29274 18814 29274 0 _0839_
rlabel viali 16692 31314 16692 31314 0 _0840_
rlabel metal2 18630 30838 18630 30838 0 _0841_
rlabel metal1 18354 29682 18354 29682 0 _0842_
rlabel metal3 17365 10404 17365 10404 0 _0843_
rlabel metal1 26358 7378 26358 7378 0 _0844_
rlabel metal1 14260 30770 14260 30770 0 _0845_
rlabel metal1 14076 31790 14076 31790 0 _0846_
rlabel metal1 14214 29614 14214 29614 0 _0847_
rlabel metal1 14398 29784 14398 29784 0 _0848_
rlabel metal1 14490 29716 14490 29716 0 _0849_
rlabel metal1 13938 29750 13938 29750 0 _0850_
rlabel metal1 13478 29648 13478 29648 0 _0851_
rlabel metal2 13570 30362 13570 30362 0 _0852_
rlabel metal1 13432 9486 13432 9486 0 _0853_
rlabel metal1 18676 9962 18676 9962 0 _0854_
rlabel metal1 29302 7378 29302 7378 0 _0855_
rlabel metal1 29118 5338 29118 5338 0 _0856_
rlabel metal1 14628 33626 14628 33626 0 _0857_
rlabel metal1 14260 34034 14260 34034 0 _0858_
rlabel metal2 19274 34085 19274 34085 0 _0859_
rlabel metal1 19688 34102 19688 34102 0 _0860_
rlabel metal1 19458 33966 19458 33966 0 _0861_
rlabel metal2 20378 33660 20378 33660 0 _0862_
rlabel metal1 20286 33524 20286 33524 0 _0863_
rlabel metal1 11592 33966 11592 33966 0 _0864_
rlabel metal1 19918 33558 19918 33558 0 _0865_
rlabel metal1 19642 32844 19642 32844 0 _0866_
rlabel via3 19067 33252 19067 33252 0 _0867_
rlabel metal1 19642 5746 19642 5746 0 _0868_
rlabel metal2 17894 7004 17894 7004 0 _0869_
rlabel metal1 18860 35734 18860 35734 0 _0870_
rlabel metal1 18998 35598 18998 35598 0 _0871_
rlabel metal2 16974 34034 16974 34034 0 _0872_
rlabel metal1 16468 34102 16468 34102 0 _0873_
rlabel metal1 16790 34170 16790 34170 0 _0874_
rlabel metal1 17112 34714 17112 34714 0 _0875_
rlabel metal2 18630 33099 18630 33099 0 _0876_
rlabel metal1 17664 33626 17664 33626 0 _0877_
rlabel metal1 18492 33082 18492 33082 0 _0878_
rlabel metal1 18906 32368 18906 32368 0 _0879_
rlabel metal3 18377 32028 18377 32028 0 _0880_
rlabel metal1 18906 5678 18906 5678 0 _0881_
rlabel metal1 20102 5338 20102 5338 0 _0882_
rlabel metal1 18860 7310 18860 7310 0 _0883_
rlabel metal1 18630 7378 18630 7378 0 _0884_
rlabel metal2 19918 9248 19918 9248 0 _0885_
rlabel metal1 22356 25874 22356 25874 0 _0886_
rlabel metal2 22218 24990 22218 24990 0 _0887_
rlabel metal1 22724 25466 22724 25466 0 _0888_
rlabel metal1 20838 26282 20838 26282 0 _0889_
rlabel metal2 22678 26180 22678 26180 0 _0890_
rlabel metal1 22770 25806 22770 25806 0 _0891_
rlabel metal2 22310 24378 22310 24378 0 _0892_
rlabel metal2 21022 25500 21022 25500 0 _0893_
rlabel metal1 21022 25126 21022 25126 0 _0894_
rlabel metal1 20930 23086 20930 23086 0 _0895_
rlabel metal1 19826 9588 19826 9588 0 _0896_
rlabel metal2 19826 25942 19826 25942 0 _0897_
rlabel metal1 18998 24378 18998 24378 0 _0898_
rlabel metal2 19182 23902 19182 23902 0 _0899_
rlabel metal1 19090 23732 19090 23732 0 _0900_
rlabel metal1 19274 23562 19274 23562 0 _0901_
rlabel metal2 18722 24004 18722 24004 0 _0902_
rlabel metal1 19136 13226 19136 13226 0 _0903_
rlabel metal1 13110 24854 13110 24854 0 _0904_
rlabel metal1 12834 24888 12834 24888 0 _0905_
rlabel metal1 17626 13158 17626 13158 0 _0906_
rlabel metal1 18998 13430 18998 13430 0 _0907_
rlabel metal2 20286 9248 20286 9248 0 _0908_
rlabel metal1 19642 7854 19642 7854 0 _0909_
rlabel metal1 20608 5678 20608 5678 0 _0910_
rlabel metal1 20056 4522 20056 4522 0 _0911_
rlabel metal1 21068 5270 21068 5270 0 _0912_
rlabel metal1 30912 5202 30912 5202 0 _0913_
rlabel metal1 23092 28186 23092 28186 0 _0914_
rlabel metal2 21850 29308 21850 29308 0 _0915_
rlabel metal1 22724 29002 22724 29002 0 _0916_
rlabel metal1 22770 29138 22770 29138 0 _0917_
rlabel metal2 23230 28492 23230 28492 0 _0918_
rlabel metal1 21781 27914 21781 27914 0 _0919_
rlabel metal1 21482 28526 21482 28526 0 _0920_
rlabel metal2 17066 10710 17066 10710 0 _0921_
rlabel metal1 26864 11186 26864 11186 0 _0922_
rlabel metal1 23874 26010 23874 26010 0 _0923_
rlabel metal1 24242 27914 24242 27914 0 _0924_
rlabel metal1 24104 28050 24104 28050 0 _0925_
rlabel metal1 23276 27370 23276 27370 0 _0926_
rlabel metal1 24012 27642 24012 27642 0 _0927_
rlabel metal1 24196 26350 24196 26350 0 _0928_
rlabel metal1 23092 15470 23092 15470 0 _0929_
rlabel viali 19923 28050 19923 28050 0 _0930_
rlabel metal1 19688 27982 19688 27982 0 _0931_
rlabel metal1 19872 27914 19872 27914 0 _0932_
rlabel metal2 21482 17051 21482 17051 0 _0933_
rlabel metal1 28980 9554 28980 9554 0 _0934_
rlabel metal2 31878 9792 31878 9792 0 _0935_
rlabel metal1 33258 8874 33258 8874 0 _0936_
rlabel metal2 31970 8670 31970 8670 0 _0937_
rlabel metal2 30314 5474 30314 5474 0 _0938_
rlabel metal1 23828 35054 23828 35054 0 _0939_
rlabel metal1 21666 35666 21666 35666 0 _0940_
rlabel metal2 23690 35326 23690 35326 0 _0941_
rlabel metal1 23552 35122 23552 35122 0 _0942_
rlabel metal1 23782 33422 23782 33422 0 _0943_
rlabel metal2 23874 33660 23874 33660 0 _0944_
rlabel metal2 23782 33932 23782 33932 0 _0945_
rlabel via2 12374 16099 12374 16099 0 _0946_
rlabel metal1 25300 12274 25300 12274 0 _0947_
rlabel metal1 24196 29478 24196 29478 0 _0948_
rlabel metal1 24794 36788 24794 36788 0 _0949_
rlabel metal2 24610 36822 24610 36822 0 _0950_
rlabel metal1 24012 37910 24012 37910 0 _0951_
rlabel metal1 24472 36686 24472 36686 0 _0952_
rlabel metal1 24334 36278 24334 36278 0 _0953_
rlabel metal1 25622 36550 25622 36550 0 _0954_
rlabel metal1 23414 16490 23414 16490 0 _0955_
rlabel metal1 21942 34544 21942 34544 0 _0956_
rlabel metal1 22678 33932 22678 33932 0 _0957_
rlabel metal3 24725 17612 24725 17612 0 _0958_
rlabel metal1 25070 16082 25070 16082 0 _0959_
rlabel metal1 25392 15878 25392 15878 0 _0960_
rlabel metal1 14398 37774 14398 37774 0 _0961_
rlabel metal1 14122 35802 14122 35802 0 _0962_
rlabel metal2 13846 37094 13846 37094 0 _0963_
rlabel metal1 13754 37910 13754 37910 0 _0964_
rlabel metal1 13800 37774 13800 37774 0 _0965_
rlabel metal2 12834 36822 12834 36822 0 _0966_
rlabel metal1 12696 36210 12696 36210 0 _0967_
rlabel metal1 12190 36346 12190 36346 0 _0968_
rlabel metal1 11868 36278 11868 36278 0 _0969_
rlabel metal1 26910 16014 26910 16014 0 _0970_
rlabel metal2 18722 31552 18722 31552 0 _0971_
rlabel metal1 18216 37230 18216 37230 0 _0972_
rlabel metal1 17158 37434 17158 37434 0 _0973_
rlabel metal1 17250 37910 17250 37910 0 _0974_
rlabel via1 17894 37315 17894 37315 0 _0975_
rlabel metal1 17940 36346 17940 36346 0 _0976_
rlabel metal1 18400 37094 18400 37094 0 _0977_
rlabel metal1 18354 16592 18354 16592 0 _0978_
rlabel metal2 16790 36244 16790 36244 0 _0979_
rlabel metal3 17917 17884 17917 17884 0 _0980_
rlabel metal2 18630 17034 18630 17034 0 _0981_
rlabel metal1 19090 16082 19090 16082 0 _0982_
rlabel metal1 30544 12818 30544 12818 0 _0983_
rlabel metal1 30544 11730 30544 11730 0 _0984_
rlabel metal1 31050 11322 31050 11322 0 _0985_
rlabel metal1 27370 16014 27370 16014 0 _0986_
rlabel metal1 26772 16082 26772 16082 0 _0987_
rlabel metal1 28474 15878 28474 15878 0 _0988_
rlabel metal1 30130 11220 30130 11220 0 _0989_
rlabel metal1 32798 18258 32798 18258 0 _0990_
rlabel metal2 33166 18972 33166 18972 0 _0991_
rlabel metal1 31372 17850 31372 17850 0 _0992_
rlabel metal1 32430 18700 32430 18700 0 _0993_
rlabel metal1 35420 19346 35420 19346 0 _0994_
rlabel metal2 36294 22678 36294 22678 0 _0995_
rlabel metal1 36018 22406 36018 22406 0 _0996_
rlabel metal2 35834 21046 35834 21046 0 _0997_
rlabel metal1 36386 23188 36386 23188 0 _0998_
rlabel metal1 35696 22678 35696 22678 0 _0999_
rlabel metal1 32522 21930 32522 21930 0 _1000_
rlabel metal1 31786 31858 31786 31858 0 _1001_
rlabel metal1 32108 30226 32108 30226 0 _1002_
rlabel metal1 33258 24752 33258 24752 0 _1003_
rlabel metal1 26082 31654 26082 31654 0 _1004_
rlabel metal1 26910 30906 26910 30906 0 _1005_
rlabel metal3 27945 37332 27945 37332 0 _1006_
rlabel metal2 33074 23902 33074 23902 0 _1007_
rlabel metal2 33350 24378 33350 24378 0 _1008_
rlabel metal1 34178 24242 34178 24242 0 _1009_
rlabel metal1 34178 24106 34178 24106 0 _1010_
rlabel via1 32798 24174 32798 24174 0 _1011_
rlabel metal1 31188 28526 31188 28526 0 _1012_
rlabel metal2 31142 26588 31142 26588 0 _1013_
rlabel metal1 31786 24344 31786 24344 0 _1014_
rlabel metal1 25714 28730 25714 28730 0 _1015_
rlabel metal1 26358 29172 26358 29172 0 _1016_
rlabel metal1 27324 37774 27324 37774 0 _1017_
rlabel metal1 31694 24140 31694 24140 0 _1018_
rlabel metal1 31947 23698 31947 23698 0 _1019_
rlabel metal1 32614 23834 32614 23834 0 _1020_
rlabel metal1 32890 23120 32890 23120 0 _1021_
rlabel metal1 32890 22066 32890 22066 0 _1022_
rlabel metal2 33166 24276 33166 24276 0 _1023_
rlabel metal2 32660 24038 32660 24038 0 _1024_
rlabel metal1 32246 21896 32246 21896 0 _1025_
rlabel metal1 30774 21114 30774 21114 0 _1026_
rlabel metal1 30452 35666 30452 35666 0 _1027_
rlabel metal1 30268 35462 30268 35462 0 _1028_
rlabel metal1 29348 20434 29348 20434 0 _1029_
rlabel metal1 25990 35700 25990 35700 0 _1030_
rlabel metal2 25530 35258 25530 35258 0 _1031_
rlabel metal1 25530 20434 25530 20434 0 _1032_
rlabel metal1 27278 19788 27278 19788 0 _1033_
rlabel metal1 29854 19890 29854 19890 0 _1034_
rlabel metal1 30038 19924 30038 19924 0 _1035_
rlabel metal1 29946 19346 29946 19346 0 _1036_
rlabel metal1 30360 20434 30360 20434 0 _1037_
rlabel metal1 30406 19788 30406 19788 0 _1038_
rlabel metal2 20746 16626 20746 16626 0 _1039_
rlabel metal1 21022 17068 21022 17068 0 _1040_
rlabel via1 20378 16558 20378 16558 0 _1041_
rlabel metal1 21114 16082 21114 16082 0 _1042_
rlabel metal1 23966 11730 23966 11730 0 _1043_
rlabel metal1 20562 14348 20562 14348 0 _1044_
rlabel metal1 20792 14450 20792 14450 0 _1045_
rlabel metal2 19734 13702 19734 13702 0 _1046_
rlabel metal2 21114 13668 21114 13668 0 _1047_
rlabel metal2 22402 12852 22402 12852 0 _1048_
rlabel metal1 32982 8908 32982 8908 0 _1049_
rlabel metal1 31096 20434 31096 20434 0 _1050_
rlabel metal1 30682 19924 30682 19924 0 _1051_
rlabel metal2 35282 21828 35282 21828 0 _1052_
rlabel metal1 34638 19346 34638 19346 0 _1053_
rlabel metal1 34960 18598 34960 18598 0 _1054_
rlabel metal1 32338 17850 32338 17850 0 _1055_
rlabel metal2 29026 8398 29026 8398 0 _1056_
rlabel metal1 25622 6698 25622 6698 0 _1057_
rlabel metal1 21206 6732 21206 6732 0 _1058_
rlabel metal2 21666 10625 21666 10625 0 _1059_
rlabel metal1 25990 5202 25990 5202 0 _1060_
rlabel metal1 27094 7514 27094 7514 0 _1061_
rlabel metal1 25990 5134 25990 5134 0 _1062_
rlabel metal1 28290 8466 28290 8466 0 _1063_
rlabel metal1 29578 8976 29578 8976 0 _1064_
rlabel metal2 29762 10642 29762 10642 0 _1065_
rlabel metal1 25806 14960 25806 14960 0 _1066_
rlabel metal1 25668 13294 25668 13294 0 _1067_
rlabel metal1 26358 15470 26358 15470 0 _1068_
rlabel metal1 31786 14484 31786 14484 0 _1069_
rlabel metal1 27324 13294 27324 13294 0 _1070_
rlabel metal1 27416 11118 27416 11118 0 _1071_
rlabel metal1 27002 9520 27002 9520 0 _1072_
rlabel metal1 27186 11696 27186 11696 0 _1073_
rlabel metal1 26680 12750 26680 12750 0 _1074_
rlabel metal1 26542 13974 26542 13974 0 _1075_
rlabel metal1 26818 12852 26818 12852 0 _1076_
rlabel metal1 26082 12954 26082 12954 0 _1077_
rlabel metal1 27416 12682 27416 12682 0 _1078_
rlabel metal2 32614 17986 32614 17986 0 _1079_
rlabel metal1 33534 18394 33534 18394 0 _1080_
rlabel metal1 34454 19380 34454 19380 0 _1081_
rlabel metal1 35328 19142 35328 19142 0 _1082_
rlabel viali 35926 23086 35926 23086 0 _1083_
rlabel metal1 36064 22066 36064 22066 0 _1084_
rlabel metal1 33764 21998 33764 21998 0 _1085_
rlabel metal1 33258 24140 33258 24140 0 _1086_
rlabel metal1 33442 22066 33442 22066 0 _1087_
rlabel metal1 31326 21998 31326 21998 0 _1088_
rlabel metal2 29670 20842 29670 20842 0 _1089_
rlabel metal1 30636 20230 30636 20230 0 _1090_
rlabel metal1 22448 14994 22448 14994 0 _1091_
rlabel metal1 33672 21522 33672 21522 0 _1092_
rlabel metal1 31418 14450 31418 14450 0 _1093_
rlabel metal1 26358 19822 26358 19822 0 _1094_
rlabel metal1 30130 16116 30130 16116 0 _1095_
rlabel metal1 30820 16218 30820 16218 0 _1096_
rlabel metal1 31694 15504 31694 15504 0 _1097_
rlabel metal1 32798 15538 32798 15538 0 _1098_
rlabel metal1 29854 16014 29854 16014 0 _1099_
rlabel metal1 32798 13872 32798 13872 0 _1100_
rlabel metal1 32706 15470 32706 15470 0 _1101_
rlabel metal2 33258 13702 33258 13702 0 _1102_
rlabel metal1 33166 12886 33166 12886 0 _1103_
rlabel metal1 30866 5542 30866 5542 0 _1104_
rlabel metal1 32614 6256 32614 6256 0 _1105_
rlabel metal2 26358 4318 26358 4318 0 _1106_
rlabel metal2 23322 4794 23322 4794 0 _1107_
rlabel metal1 20010 6290 20010 6290 0 _1108_
rlabel metal1 20240 10030 20240 10030 0 _1109_
rlabel metal1 19550 6290 19550 6290 0 _1110_
rlabel metal1 23230 4658 23230 4658 0 _1111_
rlabel metal1 26174 4556 26174 4556 0 _1112_
rlabel metal1 27048 5134 27048 5134 0 _1113_
rlabel metal1 32338 5644 32338 5644 0 _1114_
rlabel metal2 32154 5508 32154 5508 0 _1115_
rlabel metal1 32384 6290 32384 6290 0 _1116_
rlabel metal2 32614 7582 32614 7582 0 _1117_
rlabel metal1 32752 8942 32752 8942 0 _1118_
rlabel metal1 33488 12750 33488 12750 0 _1119_
rlabel metal1 33442 15538 33442 15538 0 _1120_
rlabel metal1 33028 15402 33028 15402 0 _1121_
rlabel metal2 21390 12954 21390 12954 0 _1122_
rlabel metal2 20470 11594 20470 11594 0 _1123_
rlabel metal1 32706 15674 32706 15674 0 _1124_
rlabel metal1 32292 15674 32292 15674 0 _1125_
rlabel metal2 32614 15232 32614 15232 0 _1126_
rlabel metal2 30130 10438 30130 10438 0 _1127_
rlabel metal1 29762 13498 29762 13498 0 _1128_
rlabel metal1 29072 13498 29072 13498 0 _1129_
rlabel metal2 28566 13498 28566 13498 0 _1130_
rlabel metal1 32338 12784 32338 12784 0 _1131_
rlabel metal1 32706 10642 32706 10642 0 _1132_
rlabel metal1 32085 9486 32085 9486 0 _1133_
rlabel metal1 32522 9418 32522 9418 0 _1134_
rlabel metal1 29992 8942 29992 8942 0 _1135_
rlabel metal2 30406 8364 30406 8364 0 _1136_
rlabel metal1 23000 6290 23000 6290 0 _1137_
rlabel metal1 19780 7446 19780 7446 0 _1138_
rlabel metal1 21758 7888 21758 7888 0 _1139_
rlabel via1 21030 10710 21030 10710 0 _1140_
rlabel metal2 21666 10234 21666 10234 0 _1141_
rlabel metal2 22678 7922 22678 7922 0 _1142_
rlabel metal1 27508 6222 27508 6222 0 _1143_
rlabel metal1 26542 5270 26542 5270 0 _1144_
rlabel metal2 27646 5712 27646 5712 0 _1145_
rlabel metal1 27922 6800 27922 6800 0 _1146_
rlabel metal1 31786 12818 31786 12818 0 _1147_
rlabel metal1 29762 13328 29762 13328 0 _1148_
rlabel metal1 29394 12818 29394 12818 0 _1149_
rlabel metal2 22310 16388 22310 16388 0 _1150_
rlabel metal1 21528 12138 21528 12138 0 _1151_
rlabel metal1 28152 13498 28152 13498 0 _1152_
rlabel metal1 28566 15470 28566 15470 0 _1153_
rlabel metal1 32568 11118 32568 11118 0 _1154_
rlabel metal1 30682 14382 30682 14382 0 _1155_
rlabel metal1 30682 14858 30682 14858 0 _1156_
rlabel metal1 27876 15538 27876 15538 0 _1157_
rlabel via1 27370 15130 27370 15130 0 _1158_
rlabel metal2 21850 13362 21850 13362 0 _1159_
rlabel metal2 24150 13600 24150 13600 0 _1160_
rlabel metal1 27232 7174 27232 7174 0 _1161_
rlabel metal2 22862 14144 22862 14144 0 _1162_
rlabel metal1 21206 13192 21206 13192 0 _1163_
rlabel metal1 23414 13430 23414 13430 0 _1164_
rlabel metal1 24702 12784 24702 12784 0 _1165_
rlabel metal1 32614 13736 32614 13736 0 _1166_
rlabel metal1 25898 13974 25898 13974 0 _1167_
rlabel metal1 26174 13362 26174 13362 0 _1168_
rlabel metal1 25990 13940 25990 13940 0 _1169_
rlabel metal1 24886 13940 24886 13940 0 _1170_
rlabel metal1 21712 12954 21712 12954 0 _1171_
rlabel metal2 21574 13022 21574 13022 0 _1172_
rlabel metal1 23782 12342 23782 12342 0 _1173_
rlabel via1 26450 11662 26450 11662 0 _1174_
rlabel metal1 26082 10982 26082 10982 0 _1175_
rlabel metal2 25254 12580 25254 12580 0 _1176_
rlabel metal1 24380 12750 24380 12750 0 _1177_
rlabel metal1 24840 12954 24840 12954 0 _1178_
rlabel metal1 25438 13770 25438 13770 0 _1179_
rlabel metal1 28014 14824 28014 14824 0 _1180_
rlabel metal1 28290 14960 28290 14960 0 _1181_
rlabel metal1 14398 20944 14398 20944 0 _1182_
rlabel metal1 25300 19890 25300 19890 0 _1183_
rlabel metal1 33074 36006 33074 36006 0 _1184_
rlabel metal2 20378 20587 20378 20587 0 _1185_
rlabel viali 21116 20434 21116 20434 0 _1186_
rlabel metal1 21027 20944 21027 20944 0 _1187_
rlabel metal1 23414 21488 23414 21488 0 _1188_
rlabel metal1 19918 19482 19918 19482 0 _1189_
rlabel metal1 20516 20026 20516 20026 0 _1190_
rlabel metal2 23138 21182 23138 21182 0 _1191_
rlabel metal1 25254 23018 25254 23018 0 _1192_
rlabel metal1 22126 21998 22126 21998 0 _1193_
rlabel metal1 14904 15062 14904 15062 0 _1194_
rlabel metal1 15134 14926 15134 14926 0 _1195_
rlabel metal1 14858 14892 14858 14892 0 _1196_
rlabel metal1 16330 16490 16330 16490 0 _1197_
rlabel viali 15686 15467 15686 15467 0 _1198_
rlabel metal1 14214 15504 14214 15504 0 _1199_
rlabel metal1 14858 15674 14858 15674 0 _1200_
rlabel metal1 23230 21420 23230 21420 0 _1201_
rlabel metal2 24058 22338 24058 22338 0 _1202_
rlabel metal1 34822 24650 34822 24650 0 _1203_
rlabel metal1 33856 33626 33856 33626 0 _1204_
rlabel metal2 32890 13124 32890 13124 0 _1205_
rlabel metal1 32798 13498 32798 13498 0 _1206_
rlabel metal1 29578 12750 29578 12750 0 _1207_
rlabel metal1 32124 12886 32124 12886 0 _1208_
rlabel metal2 31878 13328 31878 13328 0 _1209_
rlabel metal1 25162 13226 25162 13226 0 _1210_
rlabel metal1 30636 14314 30636 14314 0 _1211_
rlabel metal1 30728 14246 30728 14246 0 _1212_
rlabel metal1 24196 8466 24196 8466 0 _1213_
rlabel metal2 24564 12852 24564 12852 0 _1214_
rlabel metal1 25990 13328 25990 13328 0 _1215_
rlabel metal1 27002 13328 27002 13328 0 _1216_
rlabel metal1 26864 12410 26864 12410 0 _1217_
rlabel metal1 27646 13498 27646 13498 0 _1218_
rlabel metal1 31464 13906 31464 13906 0 _1219_
rlabel metal1 31464 14042 31464 14042 0 _1220_
rlabel metal2 9890 19346 9890 19346 0 _1221_
rlabel metal1 30505 21998 30505 21998 0 _1222_
rlabel metal1 33626 17646 33626 17646 0 _1223_
rlabel metal2 5750 21335 5750 21335 0 _1224_
rlabel metal1 26910 21114 26910 21114 0 _1225_
rlabel metal2 26634 33286 26634 33286 0 _1226_
rlabel metal1 31832 8058 31832 8058 0 _1227_
rlabel metal1 31602 9452 31602 9452 0 _1228_
rlabel metal2 32890 10285 32890 10285 0 _1229_
rlabel metal1 26910 11084 26910 11084 0 _1230_
rlabel metal1 27186 10676 27186 10676 0 _1231_
rlabel metal1 26910 10642 26910 10642 0 _1232_
rlabel metal1 30130 10064 30130 10064 0 _1233_
rlabel metal1 30958 9554 30958 9554 0 _1234_
rlabel metal1 33626 9690 33626 9690 0 _1235_
rlabel metal1 28106 10030 28106 10030 0 _1236_
rlabel metal1 32936 6834 32936 6834 0 _1237_
rlabel metal1 30774 9112 30774 9112 0 _1238_
rlabel metal1 9430 21488 9430 21488 0 _1239_
rlabel metal2 33258 23052 33258 23052 0 _1240_
rlabel metal1 32016 21998 32016 21998 0 _1241_
rlabel metal1 32384 22746 32384 22746 0 _1242_
rlabel metal1 32292 22542 32292 22542 0 _1243_
rlabel metal1 32062 22134 32062 22134 0 _1244_
rlabel metal2 32614 21828 32614 21828 0 _1245_
rlabel metal1 13018 22610 13018 22610 0 _1246_
rlabel metal2 28520 30566 28520 30566 0 _1247_
rlabel metal1 29900 30906 29900 30906 0 _1248_
rlabel metal1 31878 7412 31878 7412 0 _1249_
rlabel metal2 30314 4794 30314 4794 0 _1250_
rlabel metal1 30268 4794 30268 4794 0 _1251_
rlabel metal1 30452 6766 30452 6766 0 _1252_
rlabel metal1 21942 7786 21942 7786 0 _1253_
rlabel metal1 23345 10710 23345 10710 0 _1254_
rlabel metal1 22218 11152 22218 11152 0 _1255_
rlabel metal1 24656 8602 24656 8602 0 _1256_
rlabel metal1 27784 8874 27784 8874 0 _1257_
rlabel via1 26818 8925 26818 8925 0 _1258_
rlabel metal1 28382 8908 28382 8908 0 _1259_
rlabel metal1 27462 9486 27462 9486 0 _1260_
rlabel metal1 28152 8942 28152 8942 0 _1261_
rlabel metal1 29394 6766 29394 6766 0 _1262_
rlabel metal1 31004 6902 31004 6902 0 _1263_
rlabel metal1 31464 6970 31464 6970 0 _1264_
rlabel metal2 21022 20587 21022 20587 0 _1265_
rlabel metal1 34362 21522 34362 21522 0 _1266_
rlabel metal1 33534 21556 33534 21556 0 _1267_
rlabel metal2 33258 20842 33258 20842 0 _1268_
rlabel metal1 33074 24616 33074 24616 0 _1269_
rlabel metal1 34316 24922 34316 24922 0 _1270_
rlabel metal1 26726 4522 26726 4522 0 _1271_
rlabel metal1 27600 4794 27600 4794 0 _1272_
rlabel metal1 28106 5066 28106 5066 0 _1273_
rlabel metal2 28014 6596 28014 6596 0 _1274_
rlabel metal1 8418 15470 8418 15470 0 clk
rlabel metal1 31280 29614 31280 29614 0 clknet_0__0514_
rlabel metal1 17894 30566 17894 30566 0 clknet_0__0515_
rlabel metal2 20010 31790 20010 31790 0 clknet_0__0516_
rlabel metal2 19550 30141 19550 30141 0 clknet_0__0517_
rlabel metal1 9522 18360 9522 18360 0 clknet_0_clk
rlabel metal1 35098 29172 35098 29172 0 clknet_1_0__leaf__0514_
rlabel metal1 10534 23120 10534 23120 0 clknet_1_0__leaf__0515_
rlabel metal1 4738 34000 4738 34000 0 clknet_1_0__leaf__0516_
rlabel metal1 9292 36142 9292 36142 0 clknet_1_0__leaf__0517_
rlabel metal1 33948 32878 33948 32878 0 clknet_1_1__leaf__0514_
rlabel metal3 20263 35972 20263 35972 0 clknet_1_1__leaf__0515_
rlabel metal1 32798 35666 32798 35666 0 clknet_1_1__leaf__0516_
rlabel metal1 29578 38420 29578 38420 0 clknet_1_1__leaf__0517_
rlabel metal1 2622 7446 2622 7446 0 clknet_2_0__leaf_clk
rlabel metal1 15640 6834 15640 6834 0 clknet_2_1__leaf_clk
rlabel metal1 1426 19414 1426 19414 0 clknet_2_2__leaf_clk
rlabel metal1 15042 25874 15042 25874 0 clknet_2_3__leaf_clk
rlabel metal1 38134 8942 38134 8942 0 cs
rlabel metal3 820 11628 820 11628 0 gpi[0]
rlabel metal3 1096 6868 1096 6868 0 gpi[1]
rlabel metal1 31096 38998 31096 38998 0 gpi[23]
rlabel metal2 10994 1554 10994 1554 0 gpi[2]
rlabel metal2 8418 1027 8418 1027 0 gpi[3]
rlabel metal1 15640 38998 15640 38998 0 gpi[4]
rlabel metal1 37444 38930 37444 38930 0 gpi[5]
rlabel metal2 37398 1027 37398 1027 0 gpi[6]
rlabel metal2 20102 39899 20102 39899 0 gpi[7]
rlabel metal1 17618 39066 17618 39066 0 gpo[0]
rlabel metal3 820 4148 820 4148 0 gpo[10]
rlabel metal2 37950 10999 37950 10999 0 gpo[11]
rlabel metal3 820 8908 820 8908 0 gpo[12]
rlabel metal2 37858 15793 37858 15793 0 gpo[13]
rlabel metal1 782 39066 782 39066 0 gpo[14]
rlabel metal1 26818 39066 26818 39066 0 gpo[15]
rlabel metal2 17434 1520 17434 1520 0 gpo[16]
rlabel metal2 46 1554 46 1554 0 gpo[17]
rlabel metal3 820 25228 820 25228 0 gpo[18]
rlabel metal2 21942 39960 21942 39960 0 gpo[19]
rlabel metal3 820 15708 820 15708 0 gpo[1]
rlabel metal1 37904 38522 37904 38522 0 gpo[20]
rlabel metal2 13202 39967 13202 39967 0 gpo[21]
rlabel metal2 3910 959 3910 959 0 gpo[22]
rlabel metal2 1978 959 1978 959 0 gpo[23]
rlabel metal2 37858 36941 37858 36941 0 gpo[24]
rlabel metal3 820 18428 820 18428 0 gpo[25]
rlabel metal2 14858 959 14858 959 0 gpo[26]
rlabel metal1 37904 34510 37904 34510 0 gpo[27]
rlabel metal3 37958 1428 37958 1428 0 gpo[28]
rlabel metal1 9200 39066 9200 39066 0 gpo[29]
rlabel metal1 38134 20774 38134 20774 0 gpo[2]
rlabel metal2 6486 959 6486 959 0 gpo[30]
rlabel metal2 12926 1520 12926 1520 0 gpo[31]
rlabel metal3 751 20468 751 20468 0 gpo[32]
rlabel via2 37858 22491 37858 22491 0 gpo[33]
rlabel metal2 19366 959 19366 959 0 gpo[3]
rlabel metal1 35604 39066 35604 39066 0 gpo[4]
rlabel metal2 33166 39423 33166 39423 0 gpo[5]
rlabel metal2 4922 39967 4922 39967 0 gpo[6]
rlabel metal1 11362 39066 11362 39066 0 gpo[7]
rlabel metal2 26450 1520 26450 1520 0 gpo[8]
rlabel metal3 1096 13668 1096 13668 0 gpo[9]
rlabel metal1 36892 18734 36892 18734 0 net1
rlabel metal1 14168 20910 14168 20910 0 net10
rlabel metal1 4922 33966 4922 33966 0 net100
rlabel metal1 13202 38318 13202 38318 0 net101
rlabel metal1 21758 38318 21758 38318 0 net102
rlabel metal1 25714 27438 25714 27438 0 net103
rlabel metal1 32752 35122 32752 35122 0 net104
rlabel metal1 33442 26996 33442 26996 0 net105
rlabel metal1 34454 31348 34454 31348 0 net106
rlabel metal1 31832 28186 31832 28186 0 net107
rlabel metal1 27692 32538 27692 32538 0 net108
rlabel metal1 25254 38318 25254 38318 0 net109
rlabel metal1 9200 36822 9200 36822 0 net11
rlabel metal1 29854 37230 29854 37230 0 net110
rlabel metal1 10258 24922 10258 24922 0 net111
rlabel metal2 9430 35943 9430 35943 0 net112
rlabel metal1 10166 28526 10166 28526 0 net113
rlabel metal1 9430 31790 9430 31790 0 net114
rlabel metal1 8832 29614 8832 29614 0 net115
rlabel metal1 8832 33490 8832 33490 0 net116
rlabel metal1 9246 38318 9246 38318 0 net117
rlabel metal1 19136 38318 19136 38318 0 net118
rlabel metal1 27554 26996 27554 26996 0 net119
rlabel metal1 18170 38522 18170 38522 0 net12
rlabel metal1 28658 34612 28658 34612 0 net120
rlabel metal1 29486 26996 29486 26996 0 net121
rlabel metal1 27278 29172 27278 29172 0 net122
rlabel metal1 29210 29172 29210 29172 0 net123
rlabel metal2 27738 31450 27738 31450 0 net124
rlabel metal1 27462 38386 27462 38386 0 net125
rlabel metal1 29118 37876 29118 37876 0 net126
rlabel metal1 28934 24820 28934 24820 0 net127
rlabel metal2 8878 5848 8878 5848 0 net128
rlabel metal1 11079 4794 11079 4794 0 net129
rlabel metal2 3910 6698 3910 6698 0 net13
rlabel metal1 9614 5270 9614 5270 0 net130
rlabel metal1 8740 6222 8740 6222 0 net131
rlabel metal1 12696 8058 12696 8058 0 net132
rlabel metal2 13846 6086 13846 6086 0 net133
rlabel metal1 16054 4624 16054 4624 0 net134
rlabel metal1 17250 5338 17250 5338 0 net135
rlabel metal1 7958 32946 7958 32946 0 net136
rlabel metal1 7498 29138 7498 29138 0 net137
rlabel metal1 8050 30260 8050 30260 0 net138
rlabel metal1 7866 31824 7866 31824 0 net139
rlabel via2 17526 10523 17526 10523 0 net14
rlabel metal1 9706 23086 9706 23086 0 net140
rlabel metal1 11270 5610 11270 5610 0 net141
rlabel metal1 2277 8942 2277 8942 0 net15
rlabel metal1 37674 16014 37674 16014 0 net16
rlabel metal2 1794 37405 1794 37405 0 net17
rlabel metal1 22862 17850 22862 17850 0 net18
rlabel metal1 17526 2414 17526 2414 0 net19
rlabel metal1 7958 14892 7958 14892 0 net2
rlabel metal2 1794 2618 1794 2618 0 net20
rlabel metal1 2024 23290 2024 23290 0 net21
rlabel metal2 22862 21097 22862 21097 0 net22
rlabel metal2 1794 15946 1794 15946 0 net23
rlabel metal1 35144 38386 35144 38386 0 net24
rlabel metal1 12742 38930 12742 38930 0 net25
rlabel metal1 4600 2414 4600 2414 0 net26
rlabel metal1 2346 2414 2346 2414 0 net27
rlabel metal1 13340 21522 13340 21522 0 net28
rlabel metal1 1932 17850 1932 17850 0 net29
rlabel metal1 8602 14994 8602 14994 0 net3
rlabel metal1 14996 2414 14996 2414 0 net30
rlabel metal2 36938 34102 36938 34102 0 net31
rlabel metal1 37352 18054 37352 18054 0 net32
rlabel metal1 9016 38522 9016 38522 0 net33
rlabel metal1 37490 20842 37490 20842 0 net34
rlabel metal1 7682 2414 7682 2414 0 net35
rlabel metal1 13064 2414 13064 2414 0 net36
rlabel metal1 1840 20910 1840 20910 0 net37
rlabel metal1 37628 22610 37628 22610 0 net38
rlabel metal2 19826 2618 19826 2618 0 net39
rlabel metal1 13662 19822 13662 19822 0 net4
rlabel metal1 35282 38522 35282 38522 0 net40
rlabel metal1 32660 38522 32660 38522 0 net41
rlabel metal1 5060 38522 5060 38522 0 net42
rlabel metal2 12374 38488 12374 38488 0 net43
rlabel metal1 19366 2312 19366 2312 0 net44
rlabel metal1 1794 13872 1794 13872 0 net45
rlabel metal1 2622 23052 2622 23052 0 net46
rlabel metal1 6670 7854 6670 7854 0 net47
rlabel metal1 6509 33422 6509 33422 0 net48
rlabel metal1 32062 16558 32062 16558 0 net49
rlabel metal1 10672 2618 10672 2618 0 net5
rlabel metal1 18216 35258 18216 35258 0 net50
rlabel metal1 14628 34170 14628 34170 0 net51
rlabel metal2 19090 26469 19090 26469 0 net52
rlabel metal1 28566 25262 28566 25262 0 net53
rlabel metal1 11776 36142 11776 36142 0 net54
rlabel metal2 22218 31824 22218 31824 0 net55
rlabel metal1 20010 24208 20010 24208 0 net56
rlabel metal1 2905 12818 2905 12818 0 net57
rlabel metal1 13885 12886 13885 12886 0 net58
rlabel metal1 5711 31790 5711 31790 0 net59
rlabel metal1 8740 2618 8740 2618 0 net6
rlabel metal1 6631 33966 6631 33966 0 net60
rlabel metal1 11355 38250 11355 38250 0 net61
rlabel metal2 33718 35938 33718 35938 0 net62
rlabel metal2 22034 37672 22034 37672 0 net63
rlabel metal1 34592 32878 34592 32878 0 net64
rlabel metal1 35144 26010 35144 26010 0 net65
rlabel metal1 34914 29274 34914 29274 0 net66
rlabel metal1 34730 25330 34730 25330 0 net67
rlabel metal1 29946 31348 29946 31348 0 net68
rlabel metal1 27002 33524 27002 33524 0 net69
rlabel metal2 15594 38743 15594 38743 0 net7
rlabel metal1 34592 33966 34592 33966 0 net70
rlabel metal1 10718 23086 10718 23086 0 net71
rlabel metal1 7038 33524 7038 33524 0 net72
rlabel metal1 6670 26996 6670 26996 0 net73
rlabel metal2 4278 30362 4278 30362 0 net74
rlabel metal1 6118 28594 6118 28594 0 net75
rlabel metal1 4186 31790 4186 31790 0 net76
rlabel metal1 8694 23732 8694 23732 0 net77
rlabel metal1 4738 26350 4738 26350 0 net78
rlabel metal2 7314 24922 7314 24922 0 net79
rlabel via2 37674 38811 37674 38811 0 net8
rlabel metal1 6854 35054 6854 35054 0 net80
rlabel metal1 7682 28084 7682 28084 0 net81
rlabel metal2 7866 31450 7866 31450 0 net82
rlabel metal1 3910 29172 3910 29172 0 net83
rlabel metal1 4278 32878 4278 32878 0 net84
rlabel metal1 8832 37230 8832 37230 0 net85
rlabel metal1 20378 37230 20378 37230 0 net86
rlabel metal1 25622 24276 25622 24276 0 net87
rlabel metal1 30590 35054 30590 35054 0 net88
rlabel metal1 30958 26350 30958 26350 0 net89
rlabel metal1 17595 2482 17595 2482 0 net9
rlabel metal2 34546 31518 34546 31518 0 net90
rlabel metal1 34822 28186 34822 28186 0 net91
rlabel metal1 31326 32538 31326 32538 0 net92
rlabel metal2 27462 36074 27462 36074 0 net93
rlabel metal1 32338 36788 32338 36788 0 net94
rlabel metal2 8694 26010 8694 26010 0 net95
rlabel metal1 5934 36142 5934 36142 0 net96
rlabel metal1 9706 27438 9706 27438 0 net97
rlabel metal1 5842 30702 5842 30702 0 net98
rlabel metal1 4094 28084 4094 28084 0 net99
rlabel metal3 820 36788 820 36788 0 nrst
rlabel metal1 38134 18054 38134 18054 0 store_en
<< properties >>
string FIXED_BBOX 0 0 39418 41562
<< end >>
