VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO stopwatch
  CLASS BLOCK ;
  FOREIGN stopwatch ;
  ORIGIN 0.000 0.000 ;
  SIZE 152.905 BY 163.625 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 25.725 10.640 27.325 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.140 10.640 62.740 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.555 10.640 98.155 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 131.970 10.640 133.570 152.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 31.060 147.440 32.660 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 66.420 147.440 68.020 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 101.780 147.440 103.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 137.140 147.440 138.740 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.425 10.640 24.025 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.840 10.640 59.440 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.255 10.640 94.855 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.670 10.640 130.270 152.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 27.760 147.440 29.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 63.120 147.440 64.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 98.480 147.440 100.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 133.840 147.440 135.440 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END clk
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 159.625 145.270 163.625 ;
    END
  END nrst
  PIN out_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END out_0[0]
  PIN out_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.390 159.625 48.670 163.625 ;
    END
  END out_0[1]
  PIN out_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END out_0[2]
  PIN out_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 148.905 54.440 152.905 55.040 ;
    END
  END out_0[3]
  PIN out_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.030 159.625 87.310 163.625 ;
    END
  END out_0[4]
  PIN out_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END out_0[5]
  PIN out_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.905 91.840 152.905 92.440 ;
    END
  END out_0[6]
  PIN out_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END out_1[0]
  PIN out_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.905 112.240 152.905 112.840 ;
    END
  END out_1[1]
  PIN out_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END out_1[2]
  PIN out_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END out_1[3]
  PIN out_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 106.350 159.625 106.630 163.625 ;
    END
  END out_1[4]
  PIN out_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 125.670 159.625 125.950 163.625 ;
    END
  END out_1[5]
  PIN out_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END out_1[6]
  PIN out_2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.290 159.625 32.570 163.625 ;
    END
  END out_2[0]
  PIN out_2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END out_2[1]
  PIN out_2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END out_2[2]
  PIN out_2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.905 13.640 152.905 14.240 ;
    END
  END out_2[3]
  PIN out_2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END out_2[4]
  PIN out_2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END out_2[5]
  PIN out_2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 12.970 159.625 13.250 163.625 ;
    END
  END out_2[6]
  PIN out_3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 148.905 34.040 152.905 34.640 ;
    END
  END out_3[0]
  PIN out_3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END out_3[1]
  PIN out_3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.905 132.640 152.905 133.240 ;
    END
  END out_3[2]
  PIN out_3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 148.905 153.040 152.905 153.640 ;
    END
  END out_3[3]
  PIN out_3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END out_3[4]
  PIN out_3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 159.625 67.990 163.625 ;
    END
  END out_3[5]
  PIN out_3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END out_3[6]
  PIN pb_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END pb_0
  PIN pb_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END pb_1
  PIN time_done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.905 71.440 152.905 72.040 ;
    END
  END time_done
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 147.200 152.405 ;
      LAYER met1 ;
        RECT 0.070 10.640 148.510 152.560 ;
      LAYER met2 ;
        RECT 0.100 159.345 12.690 160.210 ;
        RECT 13.530 159.345 32.010 160.210 ;
        RECT 32.850 159.345 48.110 160.210 ;
        RECT 48.950 159.345 67.430 160.210 ;
        RECT 68.270 159.345 86.750 160.210 ;
        RECT 87.590 159.345 106.070 160.210 ;
        RECT 106.910 159.345 125.390 160.210 ;
        RECT 126.230 159.345 144.710 160.210 ;
        RECT 145.550 159.345 148.480 160.210 ;
        RECT 0.100 4.280 148.480 159.345 ;
        RECT 0.650 3.670 15.910 4.280 ;
        RECT 16.750 3.670 35.230 4.280 ;
        RECT 36.070 3.670 54.550 4.280 ;
        RECT 55.390 3.670 73.870 4.280 ;
        RECT 74.710 3.670 93.190 4.280 ;
        RECT 94.030 3.670 109.290 4.280 ;
        RECT 110.130 3.670 128.610 4.280 ;
        RECT 129.450 3.670 147.930 4.280 ;
      LAYER met3 ;
        RECT 4.400 156.040 148.905 156.890 ;
        RECT 3.990 154.040 148.905 156.040 ;
        RECT 3.990 152.640 148.505 154.040 ;
        RECT 3.990 137.040 148.905 152.640 ;
        RECT 4.400 135.640 148.905 137.040 ;
        RECT 3.990 133.640 148.905 135.640 ;
        RECT 3.990 132.240 148.505 133.640 ;
        RECT 3.990 116.640 148.905 132.240 ;
        RECT 4.400 115.240 148.905 116.640 ;
        RECT 3.990 113.240 148.905 115.240 ;
        RECT 3.990 111.840 148.505 113.240 ;
        RECT 3.990 99.640 148.905 111.840 ;
        RECT 4.400 98.240 148.905 99.640 ;
        RECT 3.990 92.840 148.905 98.240 ;
        RECT 3.990 91.440 148.505 92.840 ;
        RECT 3.990 79.240 148.905 91.440 ;
        RECT 4.400 77.840 148.905 79.240 ;
        RECT 3.990 72.440 148.905 77.840 ;
        RECT 3.990 71.040 148.505 72.440 ;
        RECT 3.990 58.840 148.905 71.040 ;
        RECT 4.400 57.440 148.905 58.840 ;
        RECT 3.990 55.440 148.905 57.440 ;
        RECT 3.990 54.040 148.505 55.440 ;
        RECT 3.990 38.440 148.905 54.040 ;
        RECT 4.400 37.040 148.905 38.440 ;
        RECT 3.990 35.040 148.905 37.040 ;
        RECT 3.990 33.640 148.505 35.040 ;
        RECT 3.990 18.040 148.905 33.640 ;
        RECT 4.400 16.640 148.905 18.040 ;
        RECT 3.990 14.640 148.905 16.640 ;
        RECT 3.990 13.240 148.505 14.640 ;
        RECT 3.990 10.715 148.905 13.240 ;
      LAYER met4 ;
        RECT 52.735 27.375 57.440 145.345 ;
        RECT 59.840 27.375 60.740 145.345 ;
        RECT 63.140 27.375 92.855 145.345 ;
        RECT 95.255 27.375 96.155 145.345 ;
        RECT 98.555 27.375 128.270 145.345 ;
        RECT 130.670 27.375 131.570 145.345 ;
        RECT 133.970 27.375 144.145 145.345 ;
  END
END stopwatch
END LIBRARY

