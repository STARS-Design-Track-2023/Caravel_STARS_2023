magic
tech sky130A
magscale 1 2
timestamp 1694009415
<< obsli1 >>
rect 1104 2159 38272 39185
<< obsm1 >>
rect 14 2128 38442 39216
<< metal2 >>
rect 18 40762 74 41562
rect 1950 40762 2006 41562
rect 4526 40762 4582 41562
rect 6458 40762 6514 41562
rect 9034 40762 9090 41562
rect 10966 40762 11022 41562
rect 12898 40762 12954 41562
rect 15474 40762 15530 41562
rect 17406 40762 17462 41562
rect 19982 40762 20038 41562
rect 21914 40762 21970 41562
rect 24490 40762 24546 41562
rect 26422 40762 26478 41562
rect 28354 40762 28410 41562
rect 30930 40762 30986 41562
rect 32862 40762 32918 41562
rect 35438 40762 35494 41562
rect 37370 40762 37426 41562
rect 39302 40762 39358 41562
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 14830 0 14886 800
rect 17406 0 17462 800
rect 19338 0 19394 800
rect 21914 0 21970 800
rect 23846 0 23902 800
rect 26422 0 26478 800
rect 28354 0 28410 800
rect 30286 0 30342 800
rect 32862 0 32918 800
rect 34794 0 34850 800
rect 37370 0 37426 800
rect 39302 0 39358 800
<< obsm2 >>
rect 130 40706 1894 40882
rect 2062 40706 4470 40882
rect 4638 40706 6402 40882
rect 6570 40706 8978 40882
rect 9146 40706 10910 40882
rect 11078 40706 12842 40882
rect 13010 40706 15418 40882
rect 15586 40706 17350 40882
rect 17518 40706 19926 40882
rect 20094 40706 21858 40882
rect 22026 40706 24434 40882
rect 24602 40706 26366 40882
rect 26534 40706 28298 40882
rect 28466 40706 30874 40882
rect 31042 40706 32806 40882
rect 32974 40706 35382 40882
rect 35550 40706 37314 40882
rect 37482 40706 38438 40882
rect 20 856 38438 40706
rect 130 734 1894 856
rect 2062 734 3826 856
rect 3994 734 6402 856
rect 6570 734 8334 856
rect 8502 734 10910 856
rect 11078 734 12842 856
rect 13010 734 14774 856
rect 14942 734 17350 856
rect 17518 734 19282 856
rect 19450 734 21858 856
rect 22026 734 23790 856
rect 23958 734 26366 856
rect 26534 734 28298 856
rect 28466 734 30230 856
rect 30398 734 32806 856
rect 32974 734 34738 856
rect 34906 734 37314 856
rect 37482 734 38438 856
<< metal3 >>
rect 0 39448 800 39568
rect 38618 38768 39418 38888
rect 0 36728 800 36848
rect 38618 36728 39418 36848
rect 0 34688 800 34808
rect 38618 34008 39418 34128
rect 0 31968 800 32088
rect 38618 31968 39418 32088
rect 0 29928 800 30048
rect 38618 29248 39418 29368
rect 0 27208 800 27328
rect 38618 27208 39418 27328
rect 0 25168 800 25288
rect 38618 25168 39418 25288
rect 0 23128 800 23248
rect 38618 22448 39418 22568
rect 0 20408 800 20528
rect 38618 20408 39418 20528
rect 0 18368 800 18488
rect 38618 17688 39418 17808
rect 0 15648 800 15768
rect 38618 15648 39418 15768
rect 0 13608 800 13728
rect 38618 13608 39418 13728
rect 0 11568 800 11688
rect 38618 10888 39418 11008
rect 0 8848 800 8968
rect 38618 8848 39418 8968
rect 0 6808 800 6928
rect 38618 6128 39418 6248
rect 0 4088 800 4208
rect 38618 4088 39418 4208
rect 0 2048 800 2168
rect 38618 1368 39418 1488
<< obsm3 >>
rect 798 38968 38618 39201
rect 798 38688 38538 38968
rect 798 36928 38618 38688
rect 880 36648 38538 36928
rect 798 34888 38618 36648
rect 880 34608 38618 34888
rect 798 34208 38618 34608
rect 798 33928 38538 34208
rect 798 32168 38618 33928
rect 880 31888 38538 32168
rect 798 30128 38618 31888
rect 880 29848 38618 30128
rect 798 29448 38618 29848
rect 798 29168 38538 29448
rect 798 27408 38618 29168
rect 880 27128 38538 27408
rect 798 25368 38618 27128
rect 880 25088 38538 25368
rect 798 23328 38618 25088
rect 880 23048 38618 23328
rect 798 22648 38618 23048
rect 798 22368 38538 22648
rect 798 20608 38618 22368
rect 880 20328 38538 20608
rect 798 18568 38618 20328
rect 880 18288 38618 18568
rect 798 17888 38618 18288
rect 798 17608 38538 17888
rect 798 15848 38618 17608
rect 880 15568 38538 15848
rect 798 13808 38618 15568
rect 880 13528 38538 13808
rect 798 11768 38618 13528
rect 880 11488 38618 11768
rect 798 11088 38618 11488
rect 798 10808 38538 11088
rect 798 9048 38618 10808
rect 880 8768 38538 9048
rect 798 7008 38618 8768
rect 880 6728 38618 7008
rect 798 6328 38618 6728
rect 798 6048 38538 6328
rect 798 4288 38618 6048
rect 880 4008 38538 4288
rect 798 2248 38618 4008
rect 880 1968 38618 2248
rect 798 1568 38618 1968
rect 798 1395 38538 1568
<< metal4 >>
rect 4208 2128 4528 39216
rect 19568 2128 19888 39216
rect 34928 2128 35248 39216
<< obsm4 >>
rect 9075 3979 19488 38725
rect 19968 3979 29749 38725
<< labels >>
rlabel metal3 s 0 27208 800 27328 6 clk
port 1 nsew signal input
rlabel metal3 s 38618 8848 39418 8968 6 cs
port 2 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 gpi[0]
port 3 nsew signal input
rlabel metal3 s 38618 29248 39418 29368 6 gpi[10]
port 4 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 gpi[11]
port 5 nsew signal input
rlabel metal3 s 38618 13608 39418 13728 6 gpi[12]
port 6 nsew signal input
rlabel metal2 s 1950 40762 2006 41562 6 gpi[13]
port 7 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 gpi[14]
port 8 nsew signal input
rlabel metal3 s 38618 25168 39418 25288 6 gpi[15]
port 9 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 gpi[16]
port 10 nsew signal input
rlabel metal3 s 38618 4088 39418 4208 6 gpi[17]
port 11 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 gpi[18]
port 12 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 gpi[19]
port 13 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 gpi[1]
port 14 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 gpi[20]
port 15 nsew signal input
rlabel metal3 s 38618 6128 39418 6248 6 gpi[21]
port 16 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 gpi[22]
port 17 nsew signal input
rlabel metal2 s 30930 40762 30986 41562 6 gpi[23]
port 18 nsew signal input
rlabel metal2 s 28354 40762 28410 41562 6 gpi[24]
port 19 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 gpi[25]
port 20 nsew signal input
rlabel metal3 s 38618 27208 39418 27328 6 gpi[26]
port 21 nsew signal input
rlabel metal3 s 38618 31968 39418 32088 6 gpi[27]
port 22 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 gpi[28]
port 23 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 gpi[29]
port 24 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 gpi[2]
port 25 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 gpi[30]
port 26 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 gpi[31]
port 27 nsew signal input
rlabel metal2 s 24490 40762 24546 41562 6 gpi[32]
port 28 nsew signal input
rlabel metal2 s 6458 40762 6514 41562 6 gpi[33]
port 29 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 gpi[3]
port 30 nsew signal input
rlabel metal2 s 15474 40762 15530 41562 6 gpi[4]
port 31 nsew signal input
rlabel metal2 s 37370 40762 37426 41562 6 gpi[5]
port 32 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 gpi[6]
port 33 nsew signal input
rlabel metal2 s 19982 40762 20038 41562 6 gpi[7]
port 34 nsew signal input
rlabel metal2 s 39302 40762 39358 41562 6 gpi[8]
port 35 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 gpi[9]
port 36 nsew signal input
rlabel metal2 s 17406 40762 17462 41562 6 gpo[0]
port 37 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 gpo[10]
port 38 nsew signal output
rlabel metal3 s 38618 10888 39418 11008 6 gpo[11]
port 39 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 gpo[12]
port 40 nsew signal output
rlabel metal3 s 38618 15648 39418 15768 6 gpo[13]
port 41 nsew signal output
rlabel metal2 s 18 40762 74 41562 6 gpo[14]
port 42 nsew signal output
rlabel metal2 s 26422 40762 26478 41562 6 gpo[15]
port 43 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 gpo[16]
port 44 nsew signal output
rlabel metal2 s 18 0 74 800 6 gpo[17]
port 45 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 gpo[18]
port 46 nsew signal output
rlabel metal2 s 21914 40762 21970 41562 6 gpo[19]
port 47 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 gpo[1]
port 48 nsew signal output
rlabel metal3 s 38618 38768 39418 38888 6 gpo[20]
port 49 nsew signal output
rlabel metal2 s 12898 40762 12954 41562 6 gpo[21]
port 50 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 gpo[22]
port 51 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 gpo[23]
port 52 nsew signal output
rlabel metal3 s 38618 36728 39418 36848 6 gpo[24]
port 53 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 gpo[25]
port 54 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 gpo[26]
port 55 nsew signal output
rlabel metal3 s 38618 34008 39418 34128 6 gpo[27]
port 56 nsew signal output
rlabel metal3 s 38618 1368 39418 1488 6 gpo[28]
port 57 nsew signal output
rlabel metal2 s 9034 40762 9090 41562 6 gpo[29]
port 58 nsew signal output
rlabel metal3 s 38618 20408 39418 20528 6 gpo[2]
port 59 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 gpo[30]
port 60 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 gpo[31]
port 61 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 gpo[32]
port 62 nsew signal output
rlabel metal3 s 38618 22448 39418 22568 6 gpo[33]
port 63 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 gpo[3]
port 64 nsew signal output
rlabel metal2 s 35438 40762 35494 41562 6 gpo[4]
port 65 nsew signal output
rlabel metal2 s 32862 40762 32918 41562 6 gpo[5]
port 66 nsew signal output
rlabel metal2 s 4526 40762 4582 41562 6 gpo[6]
port 67 nsew signal output
rlabel metal2 s 10966 40762 11022 41562 6 gpo[7]
port 68 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 gpo[8]
port 69 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 gpo[9]
port 70 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 nrst
port 71 nsew signal input
rlabel metal3 s 38618 17688 39418 17808 6 store_en
port 72 nsew signal output
rlabel metal4 s 4208 2128 4528 39216 6 vccd1
port 73 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 39216 6 vccd1
port 73 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 39216 6 vssd1
port 74 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 39418 41562
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5132556
string GDS_FILE /home/designer-25/CUP/openlane/Eighty_Twos/runs/23_09_06_07_06/results/signoff/Eighty_Twos.magic.gds
string GDS_START 1101050
<< end >>

