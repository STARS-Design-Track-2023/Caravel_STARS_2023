* NGSPICE file created from outel8227.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

.subckt outel8227 VGND VPWR clk cs dataBusIn[0] dataBusIn[1] dataBusIn[2] dataBusIn[3]
+ dataBusIn[4] dataBusIn[5] dataBusIn[6] dataBusIn[7] dataBusOut[0] dataBusOut[1]
+ dataBusOut[2] dataBusOut[3] dataBusOut[4] dataBusOut[5] dataBusOut[6] dataBusOut[7]
+ dataBusSelect gpio[0] gpio[10] gpio[11] gpio[12] gpio[13] gpio[14] gpio[15] gpio[16]
+ gpio[17] gpio[18] gpio[19] gpio[1] gpio[20] gpio[21] gpio[22] gpio[23] gpio[24]
+ gpio[25] gpio[2] gpio[3] gpio[4] gpio[5] gpio[6] gpio[7] gpio[8] gpio[9] nrst
X_3086_ clknet_4_4_0_clk _0046_ net41 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[20\]
+ sky130_fd_sc_hd__dfrtp_2
X_2037_ _0872_ _0881_ _1002_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__o21a_1
X_2106_ _1361_ _1368_ _1373_ _1378_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__and4bb_1
X_3155_ clknet_4_2_0_clk _0113_ net34 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2939_ _0285_ _0731_ _0738_ _0350_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire29 _0973_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2655_ _0459_ _0453_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__nand2_1
X_1606_ _0879_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__buf_4
X_2724_ _0451_ _1481_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__and2b_1
X_2586_ _0444_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__clkbuf_4
X_1537_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3138_ clknet_4_11_0_clk _0098_ net45 VGND VGND VPWR VPWR gpio[7] sky130_fd_sc_hd__dfrtp_4
X_3069_ clknet_4_8_0_clk _0033_ net39 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.irqGenerated
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2440_ _0315_ _0321_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__and2_1
X_2371_ _0914_ _1317_ _1275_ _1184_ _1279_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2638_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] _0456_ VGND VGND
+ VPWR VPWR _0497_ sky130_fd_sc_hd__nand2_1
X_2707_ _0557_ _0558_ _0560_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a21oi_1
X_2569_ _0837_ _0844_ _0858_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1940_ _1208_ _1211_ _1217_ _1218_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1871_ _0976_ _1073_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2423_ top8227.internalDataflow.addressLowBusModule.busInputs\[39\] _1390_ _1391_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[31\] VGND VGND VPWR VPWR
+ _0305_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2285_ net5 _1434_ _1435_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\]
+ net19 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__a221o_1
X_2354_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _1468_ _1475_
+ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ _1307_ _1333_ _1342_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__a21oi_4
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2972_ _0161_ _0721_ _0768_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1923_ _0901_ _0854_ _1033_ _1039_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__a31o_1
X_1785_ net3 _1042_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__nor2_1
X_1854_ _1023_ _1107_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2406_ _0204_ _0286_ _0287_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__a21oi_2
X_2268_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] _1468_ _1475_
+ _0149_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__a211o_1
X_2199_ _1285_ _1471_ _0972_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__o21a_1
X_2337_ _1013_ _1009_ _1096_ _1245_ _0126_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_62_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold30 top8227.internalDataflow.stackBusModule.busInputs\[32\] VGND VGND VPWR VPWR
+ net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 top8227.demux.state_machine.currentAddress\[2\] VGND VGND VPWR VPWR net91
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_5 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1570_ _0828_ _0821_ _0820_ _0851_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__or4b_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _0972_ _1288_ _1380_ _1381_ _1382_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__a2111oi_1
X_2053_ _0818_ _1325_ _0980_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__a21o_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2955_ _0355_ _0175_ _0753_ _0730_ _0731_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2886_ _1482_ top8227.internalDataflow.accRegToDB\[6\] net22 VGND VGND VPWR VPWR
+ _0698_ sky130_fd_sc_hd__mux2_1
X_1837_ _1089_ _1095_ _1100_ _1118_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__or4_1
X_1768_ _0978_ _1058_ _1051_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__and3_1
X_1906_ _1087_ _1107_ _1186_ _1031_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__a22o_1
X_1699_ _1001_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2671_ _0524_ _0526_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__or2_1
X_1622_ _0922_ _0923_ _0924_ _0926_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__or4_1
X_2740_ _1014_ _0890_ _1214_ _1006_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a22o_1
X_1553_ top8227.PSRCurrentValue\[7\] _0847_ _0855_ top8227.PSRCurrentValue\[6\] _0857_
+ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__o221a_2
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3085_ clknet_4_5_0_clk _0045_ net41 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2036_ _0815_ _0884_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__and2_1
X_2105_ _1374_ _1360_ _1375_ _1377_ _0972_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__o41ai_4
X_3154_ clknet_4_2_0_clk _0112_ net34 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2938_ _0736_ _0730_ _0722_ _0224_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__o221a_1
X_2869_ _0687_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _0444_
+ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2723_ _0554_ _0563_ _0574_ _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2585_ _0425_ _0443_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__and2_2
X_2654_ _0453_ _0465_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__and2_1
X_1605_ _0819_ _0906_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__a21o_1
X_1536_ top8227.demux.state_machine.currentInstruction\[0\] top8227.demux.state_machine.currentInstruction\[3\]
+ top8227.demux.state_machine.currentInstruction\[2\] _0828_ VGND VGND VPWR VPWR _0841_
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3137_ clknet_4_7_0_clk _0097_ net42 VGND VGND VPWR VPWR gpio[6] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2019_ _1254_ _1291_ _1003_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__o21a_1
X_3068_ clknet_4_8_0_clk _0032_ net38 VGND VGND VPWR VPWR top8227.demux.nmi sky130_fd_sc_hd__dfrtp_4
XFILLER_0_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2370_ _0250_ _0251_ top8227.PSRCurrentValue\[0\] VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2706_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] _0457_ _0559_
+ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2637_ _0487_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__nand2_1
X_2568_ _0903_ _1346_ _0364_ _0426_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__a31o_1
X_1519_ top8227.demux.state_machine.currentInstruction\[5\] top8227.demux.state_machine.currentInstruction\[4\]
+ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__or2_1
X_2499_ _0916_ top8227.demux.setInterruptFlag _1096_ _0926_ _1006_ VGND VGND VPWR
+ VPWR _0379_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1870_ net2 _1024_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__nand2_1
X_2353_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] _1469_ _1476_
+ top8227.PSRCurrentValue\[0\] _0234_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2422_ _0161_ _0300_ _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__a21o_1
X_2284_ _0162_ _0163_ _0164_ _0165_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__o31a_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1999_ _1127_ _0887_ _1004_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1922_ _0934_ _1032_ _1024_ _1087_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__a22o_1
X_2971_ _0299_ _0722_ _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1853_ _0911_ _0871_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1784_ net61 _1035_ _1048_ _1069_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2336_ _1484_ _1492_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__mux2_1
X_2405_ _0195_ _0202_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2267_ net6 net25 _0148_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__a21o_1
X_2198_ _0955_ _1294_ _1289_ _1470_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__a211o_1
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold31 top8227.internalDataflow.stackBusModule.busInputs\[47\] VGND VGND VPWR VPWR
+ net81 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 top8227.internalDataflow.stackBusModule.busInputs\[35\] VGND VGND VPWR VPWR
+ net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 top8227.internalDataflow.stackBusModule.busInputs\[37\] VGND VGND VPWR VPWR
+ net92 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2052_ _0876_ _0834_ _0865_ _0883_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__a31oi_2
X_2121_ top8227.internalDataflow.accRegToDB\[6\] _1386_ _1393_ VGND VGND VPWR VPWR
+ _1394_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2885_ _0697_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
X_1905_ _0937_ _0846_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2954_ _0195_ _0202_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1698_ _0993_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1836_ _1106_ _1109_ _1112_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1767_ _1041_ _1044_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2319_ _0200_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__buf_2
XFILLER_0_67_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput10 net10 VGND VGND VPWR VPWR dataBusOut[0] sky130_fd_sc_hd__buf_2
XFILLER_0_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2670_ _0524_ _0526_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__and2_1
X_1621_ _0911_ _0925_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__nor2_1
X_1552_ top8227.PSRCurrentValue\[6\] _0849_ _0856_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__nand3_1
XFILLER_0_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3153_ clknet_4_2_0_clk _0111_ net34 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_2104_ _1249_ _1251_ _1258_ _1376_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__or4_2
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3084_ clknet_4_5_0_clk _0044_ net41 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2035_ _0877_ _0943_ _0944_ _0952_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2868_ _0684_ _0686_ _0477_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2937_ _0354_ _0194_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2799_ gpio[10] _0518_ _0628_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__mux2_1
X_1819_ _0939_ _0978_ _1072_ _1082_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2722_ _0458_ _0566_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2584_ _0427_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__nor2b_2
X_1604_ _0908_ _0901_ _0854_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__and3_1
X_2653_ _0269_ _0447_ _0448_ _0268_ _0510_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__a221o_2
X_1535_ _0826_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3136_ clknet_4_5_0_clk _0096_ net42 VGND VGND VPWR VPWR gpio[5] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3067_ clknet_4_11_0_clk _0031_ net38 VGND VGND VPWR VPWR top8227.demux.setInterruptFlag
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2018_ _0830_ _0842_ _0879_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2636_ _0488_ _0489_ _0492_ _0493_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__a311o_1
X_2705_ _0531_ _0549_ _0548_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1518_ _0822_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__clkbuf_4
X_2498_ top8227.PSRCurrentValue\[1\] _0368_ _0374_ _0378_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2567_ top8227.demux.nmi top8227.instructionLoader.interruptInjector.irqGenerated
+ net29 _0401_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__a2bb2oi_4
X_3119_ clknet_4_6_0_clk _0079_ net42 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2352_ net1 net25 _1478_ top8227.internalDataflow.accRegToDB\[0\] VGND VGND VPWR
+ VPWR _0234_ sky130_fd_sc_hd__a22o_1
X_2283_ _1245_ _1288_ _1384_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2421_ _0141_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2619_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] _0456_ VGND
+ VGND VPWR VPWR _0478_ sky130_fd_sc_hd__and2_1
X_1998_ top8227.branchForward _1270_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1921_ _0951_ _1033_ _1055_ _1164_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__a22o_1
X_1852_ _1123_ _1125_ _1129_ _1133_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2970_ _0355_ _1483_ _0298_ _0730_ _0731_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1783_ net2 _1050_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2266_ top8227.internalDataflow.accRegToDB\[5\] _1478_ _1469_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\]
+ _1476_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__a221o_1
X_2335_ _1331_ _0212_ _0208_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__o21a_2
X_2404_ _0224_ _0284_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_47_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2197_ _0949_ _1291_ _1002_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold32 top8227.negEdgeDetector.q1 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 top8227.internalDataflow.stackBusModule.busInputs\[45\] VGND VGND VPWR VPWR
+ net71 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 top8227.demux.state_machine.currentAddress\[4\] VGND VGND VPWR VPWR net60
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2120_ top8227.internalDataflow.stackBusModule.busInputs\[38\] _1380_ _1388_ top8227.internalDataflow.stackBusModule.busInputs\[46\]
+ _1392_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__a221o_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2051_ _1001_ _0887_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2884_ _0151_ top8227.internalDataflow.accRegToDB\[5\] net22 VGND VGND VPWR VPWR
+ _0697_ sky130_fd_sc_hd__mux2_1
X_1904_ _1038_ _1062_ _1085_ _1033_ _1184_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2953_ _0204_ _0286_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__o21a_1
X_1835_ _1036_ _1108_ _1114_ _1116_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__a211o_1
X_1697_ _0982_ _0986_ _0999_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1766_ _1025_ _1056_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2249_ _0128_ _0123_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__and2_1
X_2318_ _0127_ _0199_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
Xoutput11 net11 VGND VGND VPWR VPWR dataBusOut[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1551_ _0850_ _0851_ _0852_ _0853_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__and4b_2
X_1620_ _0850_ _0851_ _0852_ _0853_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__or4_4
X_3083_ clknet_4_5_0_clk _0043_ net42 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_3152_ clknet_4_3_0_clk _0110_ net36 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2103_ _1179_ _0950_ _0908_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__o21a_1
X_2034_ _1285_ _1306_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__nor2_1
X_2798_ _0630_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_2867_ _0320_ _0685_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__xnor2_1
X_1818_ _1096_ _1032_ _1062_ _1099_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2936_ _0216_ _0223_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1749_ net3 _1017_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__nand2_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2721_ _0458_ _0566_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__and2_1
X_2652_ _0263_ _0451_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2583_ _0985_ _0438_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__nand3_1
X_1534_ _0838_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1603_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__clkbuf_4
X_3135_ clknet_4_7_0_clk _0095_ net48 VGND VGND VPWR VPWR gpio[4] sky130_fd_sc_hd__dfrtp_4
X_3066_ clknet_4_6_0_clk _0030_ net48 VGND VGND VPWR VPWR top8227.negEdgeDetector.q1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2017_ _0981_ _1287_ _1288_ _1289_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__or4_1
XFILLER_0_70_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2919_ _1246_ _1376_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2635_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] _0455_ VGND VGND
+ VPWR VPWR _0494_ sky130_fd_sc_hd__and2_1
X_2704_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] _0457_ VGND
+ VGND VPWR VPWR _0558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2566_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__clkbuf_4
X_1517_ top8227.demux.state_machine.currentInstruction\[1\] top8227.demux.state_machine.currentInstruction\[0\]
+ _0820_ _0821_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__or4b_1
X_2497_ _0377_ _0361_ _0274_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3049_ clknet_4_13_0_clk _0018_ net48 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_3118_ clknet_4_7_0_clk _0078_ net43 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2420_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__inv_2
X_2351_ _0231_ _0232_ _1342_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__o21a_1
X_2282_ top8227.internalDataflow.accRegToDB\[4\] _1386_ _1384_ VGND VGND VPWR VPWR
+ _0164_ sky130_fd_sc_hd__a21bo_1
X_1997_ _0837_ _0844_ _0858_ _0957_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2618_ _0476_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2549_ _0414_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1920_ _1193_ _1194_ _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__or3_1
X_1851_ _0889_ _1034_ _1057_ _1099_ _1132_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1782_ top8227.demux.state_machine.currentAddress\[12\] _1035_ _1055_ _1062_ VGND
+ VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a22o_1
X_2403_ _0216_ _0223_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2265_ _1343_ _0145_ _0146_ _1342_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__a22o_1
X_2196_ _1460_ _1458_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__and2_2
XFILLER_0_41_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2334_ _1305_ _0215_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__nand2_2
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold22 top8227.internalDataflow.stackBusModule.busInputs\[43\] VGND VGND VPWR VPWR
+ net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 top8227.demux.state_machine.currentAddress\[11\] VGND VGND VPWR VPWR net61
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 top8227.internalDataflow.stackBusModule.busInputs\[34\] VGND VGND VPWR VPWR
+ net83 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2050_ _0902_ _0947_ _1320_ _1322_ _1317_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__o41a_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2952_ _0204_ _0286_ _0350_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__a21oi_1
X_1903_ _0915_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2883_ _0696_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1765_ net3 _1042_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__or2_2
X_1834_ _1038_ _1064_ _1115_ _1091_ _0950_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1696_ _0989_ _0992_ _0998_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__o21ai_1
X_2179_ _1146_ _0881_ _0941_ _1295_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__or4_1
X_2248_ _0129_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_4
X_2317_ top8227.internalDataflow.addressLowBusModule.busInputs\[27\] _0130_ _0132_
+ net4 _0198_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput12 net12 VGND VGND VPWR VPWR dataBusOut[2] sky130_fd_sc_hd__clkbuf_4
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1550_ _0849_ _0854_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3082_ clknet_4_5_0_clk _0042_ net41 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_2033_ _0912_ _1120_ _1001_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__o21a_1
X_2102_ _1209_ _0938_ _0993_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__o21a_1
X_3151_ clknet_4_2_0_clk _0109_ net36 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2935_ _0351_ _0727_ _0728_ _0735_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2797_ gpio[9] _0511_ _0628_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__mux2_1
X_2866_ _0472_ _0471_ _0674_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__o21a_1
X_1817_ _0979_ _1020_ _1098_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1748_ net4 _1017_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__nand2_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1679_ _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2651_ _0507_ _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__xnor2_1
X_1602_ top8227.demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__clkbuf_4
X_2720_ _0571_ _0572_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__xnor2_1
X_2582_ _1422_ _0439_ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1533_ _0828_ _0821_ _0820_ top8227.demux.state_machine.currentInstruction\[0\] VGND
+ VGND VPWR VPWR _0838_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3134_ clknet_4_4_0_clk _0094_ net43 VGND VGND VPWR VPWR gpio[3] sky130_fd_sc_hd__dfrtp_4
X_2016_ _0955_ _1013_ _1127_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__o21a_1
X_3065_ clknet_4_8_0_clk _0029_ net38 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2918_ _0351_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__nand2_1
X_2849_ _0497_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__nand2_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2634_ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] _0455_ VGND VGND
+ VPWR VPWR _0493_ sky130_fd_sc_hd__and2_1
X_2703_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] _0457_ VGND
+ VGND VPWR VPWR _0557_ sky130_fd_sc_hd__or2_1
X_1516_ top8227.demux.state_machine.currentInstruction\[2\] VGND VGND VPWR VPWR _0821_
+ sky130_fd_sc_hd__buf_2
X_2565_ _0982_ _0422_ _0423_ _1336_ _0976_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3117_ clknet_4_7_0_clk _0077_ net43 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_2496_ _0375_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3048_ clknet_4_13_0_clk _0017_ net49 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2350_ net1 _1434_ _1435_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
+ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__a22o_1
X_2281_ top8227.internalDataflow.addressLowBusModule.busInputs\[36\] _1390_ _1391_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[28\] VGND VGND VPWR VPWR
+ _0163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1996_ _1004_ _1016_ _1265_ _1266_ _1268_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2617_ _0424_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2548_ net85 _0274_ _0412_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux2_1
X_2479_ _0360_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1850_ _1020_ _1111_ _1130_ _1032_ _1131_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__a32o_1
X_1781_ _0987_ _1035_ _1052_ _1055_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a22o_1
X_2333_ _1312_ _0208_ _0214_ _1333_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__o22a_2
XFILLER_0_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2402_ _0260_ _0281_ _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__a21oi_4
X_2264_ net6 _1434_ _1435_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\]
+ net19 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__a221o_1
X_2195_ _1458_ _1467_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__nor2_2
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1979_ _1248_ _1249_ _1251_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold34 net17 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 top8227.demux.state_machine.timeState\[3\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 top8227.instructionLoader.interruptInjector.irqGenerated VGND VGND VPWR VPWR
+ net62 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1902_ _1173_ _1174_ _1178_ _1182_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__or4_1
X_2951_ _1261_ _0726_ _0748_ _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__or4b_1
XFILLER_0_52_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2882_ _0174_ top8227.internalDataflow.accRegToDB\[4\] net22 VGND VGND VPWR VPWR
+ _0696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1833_ _1097_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__inv_2
X_1764_ _1054_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2316_ top8227.internalDataflow.addressLowBusModule.busInputs\[35\] net24 _0125_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] _0126_ VGND VGND VPWR
+ VPWR _0198_ sky130_fd_sc_hd__a221o_1
X_1695_ _0993_ _0994_ _0995_ _0996_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__o221a_1
X_2247_ _0128_ _0123_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2178_ _1446_ _1447_ _1450_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__and3_1
Xoutput13 net13 VGND VGND VPWR VPWR dataBusOut[3] sky130_fd_sc_hd__buf_2
XFILLER_0_31_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3150_ clknet_4_9_0_clk _0108_ net44 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3081_ clknet_4_5_0_clk _0041_ net41 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2101_ _0891_ _0923_ _0951_ _0993_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__o31a_1
X_2032_ _1304_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__buf_2
XFILLER_0_72_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2865_ _0682_ _0683_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2934_ _0733_ _0734_ top8227.internalDataflow.addressLowBusModule.busInputs\[25\]
+ _0717_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2796_ _0629_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1678_ _0980_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1747_ net2 _1017_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__nand2_2
X_1816_ _1040_ _1018_ _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__a21oi_4
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2650_ _0480_ _0500_ _0478_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__a21oi_1
X_1601_ _0902_ _0904_ _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__or3_1
X_2581_ top8227.demux.state_machine.currentAddress\[6\] _1273_ VGND VGND VPWR VPWR
+ _0440_ sky130_fd_sc_hd__nand2_1
X_1532_ top8227.PSRCurrentValue\[0\] _0823_ _0826_ _0831_ _0836_ VGND VGND VPWR VPWR
+ _0837_ sky130_fd_sc_hd__o311a_1
XFILLER_0_22_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3133_ clknet_4_8_0_clk _0093_ net38 VGND VGND VPWR VPWR gpio[2] sky130_fd_sc_hd__dfrtp_4
X_2015_ _1096_ _1275_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__and2_1
X_3064_ clknet_4_8_0_clk _0028_ net45 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.resetDetected
+ sky130_fd_sc_hd__dfstp_1
X_2848_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] _0458_ VGND VGND
+ VPWR VPWR _0669_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2917_ _0718_ _0258_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__xor2_1
X_2779_ top8227.instructionLoader.interruptInjector.resetDetected _0986_ _0402_ top8227.demux.reset
+ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__a22o_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2702_ _0503_ _0550_ _0551_ _0556_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2633_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _0490_ _0491_
+ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__a21o_1
X_1515_ top8227.demux.state_machine.currentInstruction\[3\] VGND VGND VPWR VPWR _0820_
+ sky130_fd_sc_hd__buf_2
X_2564_ _0909_ _1270_ _1427_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__nor3_1
X_2495_ _0316_ _1494_ _0153_ _0374_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3116_ clknet_4_6_0_clk _0076_ net42 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3047_ clknet_4_13_0_clk _0016_ net49 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2280_ top8227.internalDataflow.stackBusModule.busInputs\[36\] _1380_ _1388_ top8227.internalDataflow.stackBusModule.busInputs\[44\]
+ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2616_ _0453_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1995_ _1267_ top8227.demux.state_machine.currentAddress\[12\] _0965_ VGND VGND VPWR
+ VPWR _1268_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2547_ _0413_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2478_ _1246_ _0359_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1780_ net59 _1035_ _1068_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a21bo_1
X_2332_ _1343_ _0212_ _0213_ _1342_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a22o_1
X_2401_ _0282_ _0280_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__nor2_1
X_2194_ _1460_ _1466_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__or2_1
X_2263_ _1384_ _0144_ net20 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1978_ _0908_ _1250_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__and2_2
XFILLER_0_15_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold35 net11 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 top8227.internalDataflow.addressLowBusModule.busInputs\[24\] VGND VGND VPWR
+ VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 top8227.internalDataflow.addressLowBusModule.busInputs\[30\] VGND VGND VPWR
+ VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2881_ _0695_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1832_ _1020_ _1111_ _1113_ _1091_ _0949_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__a32o_1
X_2950_ _0289_ _0291_ _0741_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__or3_1
X_1901_ _1179_ _1092_ _1055_ _1107_ _1181_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1763_ net2 _0978_ _1018_ net1 VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__and4b_1
X_1694_ _0907_ top8227.demux.state_machine.currentAddress\[5\] VGND VGND VPWR VPWR
+ _0997_ sky130_fd_sc_hd__nand2_1
X_2246_ _1506_ _0118_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__nor2_1
X_2315_ _1484_ _1492_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_1
X_2177_ _0987_ _1275_ _1449_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput14 net14 VGND VGND VPWR VPWR dataBusOut[4] sky130_fd_sc_hd__clkbuf_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3080_ clknet_4_7_0_clk _0040_ net48 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
X_2100_ _0969_ _0983_ _1372_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__or3_2
XFILLER_0_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2031_ _1284_ _0985_ _1300_ _1303_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__and4b_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2864_ _0499_ _0481_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__and2b_1
X_2795_ gpio[8] _0453_ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2933_ _0283_ _0731_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__nor2_1
X_1815_ _1022_ _1049_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1677_ top8227.demux.isAddressing net33 VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__and2_1
X_1746_ top8227.demux.state_machine.currentAddress\[6\] _1035_ _1039_ _1040_ VGND
+ VGND VPWR VPWR _0009_ sky130_fd_sc_hd__a22o_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ _0916_ _0965_ _0896_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1600_ _0883_ _0864_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__nor2_2
X_2580_ _1002_ _0421_ _1016_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__o21ai_1
X_1531_ _0832_ _0834_ _0835_ top8227.PSRCurrentValue\[7\] VGND VGND VPWR VPWR _0836_
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3132_ clknet_4_11_0_clk _0092_ net45 VGND VGND VPWR VPWR gpio[1] sky130_fd_sc_hd__dfrtp_4
X_3063_ clknet_4_9_0_clk _0027_ net45 VGND VGND VPWR VPWR top8227.freeCarry sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2014_ _1209_ _0949_ _1002_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2847_ _0485_ _0472_ _0496_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2778_ _0613_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
X_2916_ _0259_ _0249_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__or2b_1
X_1729_ net5 VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__buf_2
XFILLER_0_13_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2701_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] _0445_ _0555_
+ _0477_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__a22o_1
X_2632_ _0442_ _0426_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\]
+ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1514_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2563_ _1016_ top8227.demux.state_machine.currentAddress\[6\] _1428_ _0421_ _1267_
+ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__o221ai_1
X_2494_ _0176_ _0196_ _0217_ _0358_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__or4_1
X_3115_ clknet_4_7_0_clk _0075_ net42 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_3046_ clknet_4_13_0_clk _0015_ net48 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1994_ top8227.demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2615_ _0459_ _0465_ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2546_ net10 _0358_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2477_ _0886_ _1184_ _1014_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3029_ top8227.PSRCurrentValue\[7\] _0316_ _0812_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2400_ _1305_ _0271_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2331_ net3 _1434_ _1435_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\]
+ net19 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__a221o_1
X_2262_ top8227.internalDataflow.accRegToDB\[5\] _1386_ _0143_ VGND VGND VPWR VPWR
+ _0144_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2193_ _0969_ _0983_ _1465_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__or3b_1
X_1977_ _0839_ _0846_ _0928_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2529_ _0401_ _0986_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__nor2_1
Xhold25 top8227.internalDataflow.addressHighBusModule.busInputs\[16\] VGND VGND VPWR
+ VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 top8227.pulse_slower.currentEnableState\[0\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 net15 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2880_ _0193_ top8227.internalDataflow.accRegToDB\[3\] _0691_ VGND VGND VPWR VPWR
+ _0695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1831_ _0978_ _1057_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1900_ _1180_ _1091_ _1087_ _1164_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1693_ _0907_ _0818_ _0814_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__or3b_2
X_1762_ net54 _1035_ _1053_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a21o_1
X_2314_ _1493_ _0190_ _0186_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__o21a_2
X_2245_ _1439_ _0126_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__and2_1
X_2176_ _0993_ _1448_ _1265_ top8227.demux.state_machine.currentAddress\[6\] VGND
+ VGND VPWR VPWR _1449_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput15 net15 VGND VGND VPWR VPWR dataBusOut[5] sky130_fd_sc_hd__clkbuf_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ _0987_ _1262_ _1302_ _1004_ _1078_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2932_ _0729_ _0730_ _0731_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2863_ _0482_ _0679_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__nor2_1
X_1814_ _0896_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__buf_4
X_2794_ _0614_ _0616_ _0986_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__o211a_4
XFILLER_0_40_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1745_ net6 VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__buf_2
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1676_ _0978_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__buf_4
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2159_ _0981_ _1306_ _1427_ _1431_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__o31a_1
X_2228_ _1264_ _1429_ _1499_ _1500_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1530_ top8227.demux.state_machine.currentInstruction\[4\] VGND VGND VPWR VPWR _0835_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3131_ clknet_4_7_0_clk _0091_ net48 VGND VGND VPWR VPWR gpio[0] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2013_ _0923_ _0950_ _1003_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__o21a_1
X_3062_ clknet_4_9_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
+ net38 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2915_ _0342_ net32 _0716_ _1491_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__a31o_4
XFILLER_0_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2846_ _0159_ _0666_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__xnor2_1
X_2777_ net81 _0314_ _0605_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__mux2_1
X_1728_ net6 _1023_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__and2_2
X_1659_ _0958_ _0959_ _0961_ _0963_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__a31oi_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2700_ _0553_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__xnor2_1
X_2631_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] _0442_ _0426_
+ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__or3_1
X_2562_ _0955_ _0901_ _0854_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1513_ top8227.demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2493_ _1345_ _0373_ _1246_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__o21ai_1
X_3045_ clknet_4_13_0_clk _0014_ net48 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_3114_ clknet_4_4_0_clk _0074_ net40 VGND VGND VPWR VPWR gpio[15] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2829_ _0494_ _0488_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout50 net9 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1993_ _0987_ top8227.demux.state_machine.currentAddress\[6\] VGND VGND VPWR VPWR
+ _1266_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2614_ _0320_ _0471_ _0472_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2545_ _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2476_ _1493_ _0245_ _0237_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3028_ _1344_ _0373_ _0811_ _1247_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__o31a_1
XFILLER_0_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2192_ _1078_ _1462_ _1464_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__a21oi_2
X_2330_ _1384_ _0211_ net20 VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a21oi_2
X_2261_ top8227.internalDataflow.stackBusModule.busInputs\[37\] _1380_ _1388_ top8227.internalDataflow.stackBusModule.busInputs\[45\]
+ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1976_ _0894_ _0854_ _1084_ _0908_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2528_ net55 VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__inv_2
Xhold26 top8227.internalDataflow.addressHighBusModule.busInputs\[22\] VGND VGND VPWR
+ VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 top8227.internalDataflow.stackBusModule.busInputs\[44\] VGND VGND VPWR VPWR
+ net65 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 top8227.internalDataflow.stackBusModule.busInputs\[36\] VGND VGND VPWR VPWR
+ net87 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ _0340_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__buf_2
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1830_ _1110_ _1032_ _1087_ _1111_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1761_ _0979_ _1020_ _1052_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__and3_2
XFILLER_0_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2313_ _0194_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__inv_2
X_1692_ top8227.demux.state_machine.currentAddress\[10\] top8227.demux.state_machine.currentAddress\[4\]
+ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2244_ _0119_ _0123_ _0125_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__nor3_4
X_2175_ _1016_ _1301_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1959_ _1155_ _1159_ _1177_ _1187_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__or4_1
Xoutput16 net16 VGND VGND VPWR VPWR dataBusOut[6] sky130_fd_sc_hd__buf_2
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2931_ _0283_ _0729_ _0722_ _0216_ _0355_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__o32a_1
X_2862_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] _0445_ _0678_
+ _0477_ _0681_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__a221o_1
X_2793_ _1407_ _0617_ _0622_ _0626_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1744_ _1023_ _1036_ _1038_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__and3_1
X_1813_ _1090_ _1092_ _1038_ _1094_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__a22o_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1675_ _0976_ _0977_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__nor2_2
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2158_ _1078_ _1429_ _1430_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__or3_1
X_2227_ _1267_ _0987_ _0965_ _1448_ _1262_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__a32o_1
X_2089_ _0902_ _1131_ _1195_ _0949_ _0993_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__o41a_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3130_ clknet_4_1_0_clk _0090_ net40 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2012_ top8227.branchBackward _1270_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__and2_1
X_3061_ clknet_4_9_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
+ net39 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[3\] sky130_fd_sc_hd__dfrtp_2
X_2845_ _0472_ _0470_ _0660_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__o21a_1
X_2914_ _0353_ _0346_ _0715_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__nor3_1
X_1658_ top8227.demux.reset _0962_ _0894_ _0849_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2776_ _0612_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
X_1727_ _1021_ _1022_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__nor2_1
X_1589_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__clkbuf_4
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2561_ _0420_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
X_2630_ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] _0455_ VGND VGND
+ VPWR VPWR _0489_ sky130_fd_sc_hd__xor2_1
X_1512_ _0815_ _0816_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2492_ _0369_ _1351_ _0370_ _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__or4_2
XFILLER_0_42_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3113_ clknet_4_5_0_clk _0073_ net44 VGND VGND VPWR VPWR gpio[14] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3044_ clknet_4_15_0_clk _0013_ net48 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_2828_ _0648_ _0651_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__nand2_1
X_2759_ _0932_ _0944_ _1197_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__or3_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout40 net41 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1992_ _0957_ _0815_ _0908_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__a21o_2
XFILLER_0_42_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2613_ _0455_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2544_ _0985_ _0408_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2475_ _1261_ _0331_ _0334_ _0352_ _0356_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__o32a_2
XFILLER_0_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3027_ _1015_ _0923_ _0387_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2191_ _1226_ _1463_ _1078_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__a21oi_1
X_2260_ top8227.internalDataflow.addressLowBusModule.busInputs\[37\] _1390_ _1391_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[29\] VGND VGND VPWR VPWR
+ _0142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1975_ _1002_ _0903_ _0854_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__and3_2
XFILLER_0_43_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold38 top8227.internalDataflow.addressLowBusModule.busInputs\[20\] VGND VGND VPWR
+ VPWR net88 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold16 top8227.internalDataflow.stackBusModule.busInputs\[46\] VGND VGND VPWR VPWR
+ net66 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2458_ top8227.PSRCurrentValue\[3\] _1246_ _0250_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__and3_1
Xhold27 top8227.demux.state_machine.currentAddress\[10\] VGND VGND VPWR VPWR net77
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2527_ _0400_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
X_2389_ _1312_ _0264_ _0270_ _1333_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__o22a_2
XFILLER_0_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1760_ _1044_ _1051_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__nor2_2
X_1691_ top8227.demux.state_machine.currentAddress\[7\] top8227.demux.state_machine.currentAddress\[3\]
+ top8227.demux.state_machine.currentAddress\[11\] _0818_ VGND VGND VPWR VPWR _0994_
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_57_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2312_ _1305_ _0193_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2243_ _0124_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_4
X_2174_ _1263_ _1317_ _0971_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput17 net17 VGND VGND VPWR VPWR dataBusOut[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1889_ _0946_ _1092_ _1080_ _1087_ _1169_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1958_ _1038_ _1234_ _1213_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2861_ _0679_ _0503_ _0680_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__and3b_1
XFILLER_0_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2930_ _1246_ _1376_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__nand2_4
X_2792_ _0910_ _1410_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__or3_1
XFILLER_0_40_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1674_ top8227.instructionLoader.interruptInjector.resetDetected gpio[21] VGND VGND
+ VPWR VPWR _0977_ sky130_fd_sc_hd__nor2_1
X_1812_ _1027_ _1047_ _1093_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__a21oi_1
X_1743_ _1037_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__clkbuf_4
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _1267_ top8227.demux.state_machine.currentAddress\[12\] _1498_ VGND VGND VPWR
+ VPWR _1499_ sky130_fd_sc_hd__and3_1
X_2157_ top8227.demux.state_machine.currentAddress\[12\] _0990_ _0991_ _1262_ _1016_
+ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__a32o_1
X_2088_ top8227.pulse_slower.nextEnableState\[0\] _0974_ _1356_ _1360_ _0972_ VGND
+ VGND VPWR VPWR _1361_ sky130_fd_sc_hd__a32o_2
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3060_ clknet_4_9_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
+ net38 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2011_ _1264_ _1269_ _1271_ _1283_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2844_ net88 _0445_ _0663_ _0477_ _0665_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2913_ _0982_ _1286_ net31 _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__or4bb_1
X_1657_ top8227.demux.state_machine.timeState\[4\] _0814_ top8227.demux.state_machine.timeState\[6\]
+ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__nor3_1
X_1588_ _0821_ _0820_ _0828_ top8227.demux.state_machine.currentInstruction\[0\] VGND
+ VGND VPWR VPWR _0893_ sky130_fd_sc_hd__and4b_1
X_2775_ net66 _1482_ _0605_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1726_ net7 _1017_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__nand2_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2209_ _1442_ _1481_ _1333_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__mux2_2
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2560_ net84 _0316_ _0412_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__mux2_1
X_1511_ top8227.branchBackward top8227.branchForward VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__nor2_1
X_2491_ _1309_ _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3112_ clknet_4_1_0_clk _0072_ net40 VGND VGND VPWR VPWR gpio[13] sky130_fd_sc_hd__dfrtp_4
X_3043_ clknet_4_11_0_clk _0003_ net45 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_73_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2827_ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] _0445_ _0650_
+ _0425_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2758_ _0601_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
X_2689_ _0425_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__nor2_1
X_1709_ _1000_ _0977_ _0986_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__and3b_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout41 net44 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_4
XFILLER_0_51_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2612_ _0135_ _0159_ _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1991_ _1262_ _1263_ _1078_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2543_ _1006_ _1294_ _0882_ _1015_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2474_ _0239_ _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__nor2_1
X_3026_ top8227.demux.isAddressing _0979_ _0810_ _1010_ VGND VGND VPWR VPWR _0116_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2190_ _0988_ _0992_ _0998_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1974_ _1246_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__buf_4
XFILLER_0_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2388_ _1343_ _0268_ _0269_ _1342_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold39 top8227.internalDataflow.stackBusModule.busInputs\[39\] VGND VGND VPWR VPWR
+ net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 top8227.internalDataflow.addressLowBusModule.busInputs\[31\] VGND VGND VPWR
+ VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 top8227.demux.setInterruptFlag VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2526_ top8227.freeCarry _0357_ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux2_1
X_2457_ _0322_ _0338_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__nor2_1
X_3009_ _0801_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1690_ _0907_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__clkbuf_4
X_2311_ _1312_ _0186_ _0192_ _1333_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__o22a_2
X_2242_ _0122_ _1497_ _0118_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__and3b_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2173_ top8227.demux.state_machine.currentAddress\[12\] _1265_ VGND VGND VPWR VPWR
+ _1446_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1957_ _1051_ _1056_ _1103_ _1233_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__a31o_1
Xoutput18 net18 VGND VGND VPWR VPWR dataBusSelect sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2509_ _1006_ _0950_ _0359_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__a21oi_1
X_1888_ _0952_ _1091_ _1054_ _1103_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2860_ _0484_ _0498_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2791_ _1406_ _1399_ _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1811_ _1040_ net7 _1049_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__or3_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1673_ _0975_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1742_ _0978_ _1019_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__and2_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _0957_ _0960_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2156_ _1267_ _1428_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__and2_1
X_2087_ _1359_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2989_ _0329_ _0784_ _0334_ _0781_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__o31a_1
XFILLER_0_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2010_ _1272_ _1277_ _1280_ _1282_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__or4_1
XFILLER_0_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2912_ _1249_ _1251_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2843_ _0487_ _0495_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2774_ _0611_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
X_1725_ net8 VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__buf_4
X_1656_ _0960_ _0879_ _0864_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__or3_1
X_1587_ _0815_ _0890_ _0891_ _0819_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__a22o_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2139_ _1400_ _1411_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__and2_1
X_2208_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] _1468_ _1475_
+ _1480_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__a211o_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1510_ _0814_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__buf_2
X_2490_ _0891_ _0934_ _1327_ _1015_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__o31a_1
XFILLER_0_65_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3111_ clknet_4_5_0_clk _0071_ net44 VGND VGND VPWR VPWR gpio[12] sky130_fd_sc_hd__dfrtp_4
X_3042_ clknet_4_12_0_clk _0002_ net46 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2688_ _0536_ _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2826_ _0222_ _0649_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2757_ _0314_ top8227.internalDataflow.addressLowBusModule.busInputs\[39\] _0593_
+ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__mux2_1
X_1708_ _0976_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__buf_4
X_1639_ _0901_ _0921_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__and2_2
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout42 net43 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_4
XFILLER_0_51_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1990_ top8227.demux.state_machine.currentAddress\[10\] top8227.demux.state_machine.currentAddress\[4\]
+ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__or2_2
X_2611_ _0180_ _0427_ _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__and3_1
X_2542_ _1127_ _1274_ _1288_ _0982_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__a211o_1
X_2473_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__inv_2
X_3025_ _0809_ _0999_ top8227.demux.isAddressing VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2809_ gpio[15] _0587_ _0628_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1973_ _1245_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2525_ _0982_ _1298_ _0398_ _0986_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__o211a_1
X_2387_ net2 _1434_ _1435_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
+ _1440_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold18 top8227.internalDataflow.stackBusModule.busInputs\[42\] VGND VGND VPWR VPWR
+ net68 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 net12 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
X_2456_ _0141_ _0337_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__and2_1
X_3008_ top8227.internalDataflow.stackBusModule.busInputs\[33\] _0271_ _0799_ VGND
+ VGND VPWR VPWR _0801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2172_ _1443_ _1444_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__nor2_1
X_2310_ _1343_ _0190_ _0191_ _1342_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__a22o_1
X_2241_ _1497_ _0122_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1887_ _0884_ _1092_ _1057_ _1082_ _1167_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1956_ net4 _1093_ _1018_ _1025_ net3 VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2508_ _1246_ _0250_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nand2_1
X_2439_ _0317_ _0320_ _0139_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__mux2_1
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2790_ _1294_ _1275_ _1347_ _0433_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_25_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1741_ _1025_ _1026_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1810_ _1091_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1672_ top8227.pulse_slower.nextEnableState\[0\] _0974_ VGND VGND VPWR VPWR _0975_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _1437_ _1496_ _0972_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__o21ai_1
X_2155_ _0819_ _0991_ top8227.demux.state_machine.currentAddress\[6\] VGND VGND VPWR
+ VPWR _1428_ sky130_fd_sc_hd__o21a_1
X_2086_ _1357_ _1358_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1939_ _1124_ _1132_ _1174_ _1193_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2988_ _0325_ _0326_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2911_ _0320_ _0713_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2842_ _0496_ _0503_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2773_ net71 _0151_ _0605_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1724_ _1019_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__clkbuf_4
X_1655_ top8227.demux.state_machine.timeState\[2\] top8227.demux.state_machine.timeState\[6\]
+ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__nor2_2
X_1586_ _0874_ _0871_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__nor2_4
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2069_ _1341_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__clkbuf_4
X_2138_ _0834_ _0885_ _0883_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_48_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\] _1469_ _1476_
+ top8227.PSRCurrentValue\[6\] _1479_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__a221o_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3110_ clknet_4_7_0_clk _0070_ net42 VGND VGND VPWR VPWR gpio[11] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_50_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3041_ clknet_4_10_0_clk _0001_ net46 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2825_ _0459_ _0467_ _0460_ _0539_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1707_ top8227.demux.state_machine.timeState\[1\] VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__clkbuf_4
X_2687_ _0541_ _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__nand2_1
X_1638_ _0883_ _0925_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__nor2_2
XFILLER_0_41_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2756_ _0600_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1569_ _0873_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__buf_4
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout43 net44 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2610_ _0201_ _0468_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2541_ _1315_ _1464_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__nand2_1
X_2472_ _1249_ _0353_ _1245_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__o21a_1
X_3024_ top8227.demux.state_machine.currentAddress\[8\] top8227.demux.state_machine.currentAddress\[0\]
+ top8227.demux.state_machine.currentAddress\[2\] top8227.demux.state_machine.currentAddress\[9\]
+ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2808_ _0635_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2739_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\] _0445_ _0584_
+ _0503_ _0590_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1972_ _0972_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2524_ _0987_ _1262_ _1422_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2455_ _0161_ _0336_ _0303_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__a21o_1
X_2386_ _1384_ _0265_ _0266_ _0267_ net93 VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold19 top8227.internalDataflow.addressLowBusModule.busInputs\[29\] VGND VGND VPWR
+ VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3007_ _0800_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2171_ _0819_ _0896_ _0912_ _0815_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__a22o_1
X_2240_ _0984_ _1501_ _1505_ _0121_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1886_ _1072_ _1086_ _1093_ _1091_ _0932_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1955_ _0943_ _1034_ _1143_ _1149_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2438_ _0127_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__nand2b_4
X_2507_ _0196_ _0361_ _0385_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2369_ _0881_ _0934_ _1186_ _1004_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__o31a_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1671_ _0971_ _0968_ gpio[19] VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1740_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _0916_ _0896_ _0914_ _1013_ _1426_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__a221o_1
X_2223_ _1002_ _1009_ _1127_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__o21a_1
X_2085_ _0886_ _0932_ _1321_ _0908_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__o31a_1
X_2987_ _0741_ _0782_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1869_ _0874_ _0839_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1938_ _1100_ _1213_ _1215_ _1216_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__or4b_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2841_ _0659_ _0660_ _0662_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__o21bai_1
X_2910_ gpio[7] _0708_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__nand2_1
X_1654_ _0849_ _0894_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__nand2_1
X_2772_ _0610_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
X_1723_ net1 net2 _1018_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__o21ai_1
X_1585_ _0874_ _0823_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__nor2_2
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ net7 net25 _1478_ top8227.internalDataflow.accRegToDB\[6\] VGND VGND VPWR
+ VPWR _1479_ sky130_fd_sc_hd__a22o_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2137_ _1400_ _1151_ _0952_ _1316_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__a22o_1
X_2068_ _0972_ _1312_ _1334_ _1340_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3040_ clknet_4_10_0_clk _0012_ net47 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2824_ _0646_ _0477_ _0443_ _0647_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1706_ _1008_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
X_2686_ _0472_ _0511_ _0512_ _0518_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__nand4_1
X_1637_ _0876_ _0920_ _0826_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2755_ _1482_ top8227.internalDataflow.addressLowBusModule.busInputs\[38\] _0593_
+ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__mux2_1
X_1568_ _0835_ _0832_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__or2b_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout44 net50 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2471_ _0877_ _1151_ _1005_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__o21a_1
X_2540_ net62 _0405_ _0407_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__a21bo_1
X_3023_ _0357_ _0808_ _0396_ net57 VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2807_ gpio[14] _0578_ _0628_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2738_ _0588_ _0589_ _0425_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2669_ _0480_ _0500_ _0525_ _0506_ _0478_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__a311o_1
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1971_ gpio[16] VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiSync.in
+ sky130_fd_sc_hd__inv_2
X_2523_ net56 _0396_ _0397_ _0357_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2385_ top8227.internalDataflow.accRegToDB\[1\] _1386_ VGND VGND VPWR VPWR _0267_
+ sky130_fd_sc_hd__nand2_1
X_2454_ _0182_ _0335_ _0299_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__a21o_1
X_3006_ net80 _0238_ _0799_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__mux2_1
Xinput1 dataBusIn[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2170_ _1001_ _0889_ _0896_ _1014_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__a22o_1
X_1954_ _1231_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1885_ _0898_ _1092_ _1072_ _1099_ _1165_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2437_ top8227.internalDataflow.addressLowBusModule.busInputs\[31\] _0130_ _0132_
+ _1021_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__a221o_1
X_2506_ _0364_ _0363_ _0383_ _0384_ top8227.PSRCurrentValue\[3\] VGND VGND VPWR VPWR
+ _0385_ sky130_fd_sc_hd__a32o_1
X_2368_ _1248_ _1258_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__or2_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2299_ _0177_ _0180_ _0139_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__mux2_1
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap30 net31 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1670_ net29 VGND VGND VPWR VPWR gpio[21] sky130_fd_sc_hd__clkinv_4
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _1484_ _1492_ _1494_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2153_ _0912_ _0915_ top8227.demux.state_machine.timeState\[1\] VGND VGND VPWR VPWR
+ _1426_ sky130_fd_sc_hd__o21a_1
X_2084_ _0908_ _0884_ _0958_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1937_ _0826_ _0834_ _0979_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__or3_1
X_2986_ _0781_ _0329_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1799_ _1037_ _1057_ _1080_ _1031_ _0902_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__a32o_1
X_1868_ _1146_ _1031_ _1086_ _1147_ _1149_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2840_ _0470_ _0661_ _0459_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__o21a_1
X_2771_ net65 _0174_ _0605_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1653_ _0957_ _0874_ _0936_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__or3_1
X_1584_ _0874_ _0830_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__nor2_2
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _1017_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__clkbuf_4
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _0985_ _1465_ _1458_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__and3_2
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2136_ _1406_ _1408_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__or2_1
X_2067_ _0976_ _1336_ _1339_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2969_ _0299_ _0182_ _0335_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__nand3_1
XFILLER_0_54_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1705_ _0979_ _1000_ _1007_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__or3_1
X_2823_ _0489_ _0492_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2754_ _0599_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2685_ _0537_ _0518_ _0520_ _0540_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__or4_1
X_1636_ _0823_ _0871_ _0834_ _0879_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__a31oi_4
X_1567_ _0825_ _0871_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__nor2_4
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2119_ top8227.internalDataflow.addressLowBusModule.busInputs\[38\] _1390_ _1391_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[30\] VGND VGND VPWR VPWR
+ _1392_ sky130_fd_sc_hd__a22o_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout34 net35 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
X_3099_ clknet_4_9_0_clk _0059_ net39 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[41\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout45 net47 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2470_ _0339_ _0341_ _0323_ _0351_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__o31a_1
X_3022_ _0396_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _1021_
+ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__or3b_1
XFILLER_0_58_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2668_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] _0456_ VGND
+ VGND VPWR VPWR _0525_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2737_ _0576_ _0587_ _0585_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__or3_1
X_2806_ _0634_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2599_ _0457_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__clkbuf_4
X_1619_ _0911_ _0876_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__nor2_2
XFILLER_0_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1970_ gpio[17] VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.interruptRequest
+ sky130_fd_sc_hd__inv_2
XFILLER_0_28_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2522_ _1021_ _0868_ _0364_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\]
+ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__and4b_1
XFILLER_0_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2384_ top8227.internalDataflow.addressLowBusModule.busInputs\[33\] _1390_ _1391_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[25\] VGND VGND VPWR VPWR
+ _0266_ sky130_fd_sc_hd__a22oi_2
X_2453_ _0295_ _0288_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__or2_1
X_3005_ _0797_ _0798_ _1247_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__o21a_4
Xinput2 dataBusIn[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_4
XFILLER_0_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1953_ _1225_ _1230_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1884_ _1020_ _1130_ _1164_ _1091_ _0904_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2505_ _0364_ _0383_ _0361_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__a21oi_1
X_2298_ _0127_ _0179_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__or2_4
XFILLER_0_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2436_ top8227.internalDataflow.addressLowBusModule.busInputs\[39\] net24 _0125_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _0126_ VGND VGND VPWR
+ VPWR _0318_ sky130_fd_sc_hd__a221o_1
X_2367_ _0239_ _0244_ _0248_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap20 net21 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _1396_ _1481_ _1493_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__mux2_4
X_2152_ net28 _1419_ _1421_ _1424_ _0975_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__a311o_1
X_2083_ _1345_ _1353_ _1354_ _1338_ _1355_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__o32a_1
XFILLER_0_17_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1936_ _1072_ _1086_ _1111_ _1214_ _1032_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__a32o_1
X_2985_ _0304_ _0327_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__nand2_1
X_1867_ _1087_ _1098_ _1148_ _1030_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__a22o_1
X_1798_ _1040_ _1021_ net7 _1018_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__and4b_2
X_2419_ _1483_ _0140_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2770_ _0609_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1721_ top8227.demux.nmi top8227.instructionLoader.interruptInjector.resetDetected
+ top8227.instructionLoader.interruptInjector.irqGenerated VGND VGND VPWR VPWR _1017_
+ sky130_fd_sc_hd__nor3_4
X_1652_ top8227.demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__inv_2
X_1583_ _0882_ _0887_ _0859_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__o21a_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2135_ _1294_ _0965_ _0884_ _1400_ _1407_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__a221o_1
X_2204_ _0976_ _1460_ _1465_ _1458_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__nor4_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2066_ _1078_ _1338_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2899_ gpio[0] _0708_ _0637_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2968_ _0765_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1919_ _1195_ _1033_ _1196_ _1198_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2822_ _0489_ _0492_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__and2_1
X_1704_ _1006_ top8227.demux.state_machine.timeState\[3\] _0986_ VGND VGND VPWR VPWR
+ _1007_ sky130_fd_sc_hd__mux2_1
X_2684_ _0538_ _0539_ _0320_ _0180_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_41_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2753_ _0151_ top8227.internalDataflow.addressLowBusModule.busInputs\[37\] _0593_
+ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1566_ _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__buf_4
X_1635_ _0930_ _0935_ _0938_ _0939_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__or4b_1
XFILLER_0_39_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2049_ _0993_ _1321_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__and2_1
X_2118_ _1373_ _1378_ _1361_ _1368_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__and4_4
X_3098_ clknet_4_3_0_clk _0058_ net35 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout35 net37 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
Xfanout46 net47 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3021_ _0807_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2805_ gpio[13] _0566_ _0628_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2667_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] _0457_ VGND
+ VGND VPWR VPWR _0524_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2736_ _0576_ _0585_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__o21ai_1
X_1618_ _0879_ _0920_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__nor2_4
XFILLER_0_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2598_ _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__buf_2
X_1549_ _0850_ _0851_ _0852_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2521_ _0868_ _0364_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2383_ top8227.internalDataflow.stackBusModule.busInputs\[41\] _1387_ _1381_ _1380_
+ top8227.internalDataflow.stackBusModule.busInputs\[33\] VGND VGND VPWR VPWR _0265_
+ sky130_fd_sc_hd__a32oi_4
X_2452_ _0332_ _0333_ _0323_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__a21o_1
Xinput3 dataBusIn[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XFILLER_0_52_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3004_ _0902_ _0949_ _1015_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2719_ _0557_ _0560_ _0558_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_14_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1952_ _1199_ _1227_ _1228_ _1229_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1883_ _1040_ _1021_ net7 _1018_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__and4_2
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2504_ _0849_ _0921_ _0904_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__a21o_1
X_2435_ _1484_ _1492_ _0316_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2297_ top8227.internalDataflow.addressLowBusModule.busInputs\[28\] _0130_ _0132_
+ net5 _0178_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__a221oi_4
X_2366_ _1484_ _0246_ _0247_ _0139_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap21 _1395_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap32 _1485_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2151_ top8227.demux.state_machine.currentAddress\[6\] _1265_ _1423_ VGND VGND VPWR
+ VPWR _1424_ sky130_fd_sc_hd__a21oi_1
X_2220_ _1331_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__clkbuf_4
X_2082_ _1313_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2984_ _0777_ _0779_ _0341_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__a21oi_1
X_1935_ _0834_ _0937_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__nor2_1
X_1866_ _0839_ _0937_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__nor2_1
X_1797_ _1079_ VGND VGND VPWR VPWR gpio[22] sky130_fd_sc_hd__inv_2
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2418_ _0182_ _0296_ _0299_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__a21o_1
X_2349_ _0230_ _1439_ _1434_ _1435_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_66_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1651_ _0927_ _0940_ _0954_ _0955_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1720_ top8227.demux.state_machine.currentAddress\[7\] VGND VGND VPWR VPWR _1016_
+ sky130_fd_sc_hd__clkbuf_4
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ _0884_ _0886_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__or2_2
X_2134_ _0931_ _0932_ _0933_ _0934_ _0818_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__o41a_1
X_2203_ _1458_ _1460_ _0984_ _1466_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__and4b_4
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2065_ _0995_ _0996_ _0992_ _1337_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2967_ _0762_ _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2898_ _0986_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__nand2_4
X_1849_ _0864_ _0937_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1918_ _1197_ _1091_ _1087_ _1103_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2821_ _0477_ _0641_ _0645_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__a21o_1
X_1703_ _1005_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__buf_4
X_2683_ _0472_ _0443_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__or2_1
X_1634_ _0903_ _0921_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2752_ _0598_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1565_ _0821_ _0820_ _0828_ _0851_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_39_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2048_ _0852_ _0853_ _0903_ _0850_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__and4b_4
X_2117_ _1389_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__buf_2
X_3097_ clknet_4_0_0_clk _0057_ net35 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout36 net37 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout47 net50 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
XFILLER_0_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3020_ net89 _0314_ _0799_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__mux2_1
X_2804_ _0633_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2597_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__buf_2
X_2666_ _0518_ _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__xor2_1
X_2735_ _0309_ _0447_ _0448_ _0308_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__a221o_1
X_1617_ _0874_ _0920_ _0921_ _0849_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1548_ _0820_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__clkbuf_2
X_3149_ clknet_4_3_0_clk _0107_ net36 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2520_ gpio[18] _1079_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__nand2_2
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2451_ _0141_ _0304_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__nand2_1
X_2382_ _1493_ _0263_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3003_ _0943_ _1121_ _1006_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__o21a_1
Xinput4 dataBusIn[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2718_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\] _0458_ VGND
+ VGND VPWR VPWR _0571_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2649_ _0505_ _0506_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1882_ _1163_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1951_ _1038_ _1072_ _1085_ _1034_ _0926_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2434_ _0308_ _0313_ _1493_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__mux2_2
X_2365_ _1493_ _0245_ _1492_ _0237_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2503_ _0217_ _0361_ _0382_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
+ sky130_fd_sc_hd__a21o_1
X_2296_ top8227.internalDataflow.addressLowBusModule.busInputs\[36\] net24 _0125_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] _0126_ VGND VGND VPWR
+ VPWR _0178_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap22 _0691_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2150_ _1001_ _1016_ _1422_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__a21bo_1
X_2081_ _0814_ _0868_ _1335_ _1326_ _1328_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__a311o_1
XFILLER_0_33_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2983_ _0303_ _0161_ _0336_ _0778_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__a31o_1
X_1934_ _1212_ _1091_ net26 _1107_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__a22o_1
X_1796_ _1078_ _0968_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__and2_2
XFILLER_0_24_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1865_ _1049_ _1073_ _1094_ _1139_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__nor4_1
X_2348_ _1245_ _1438_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__nand2_1
X_2417_ _0297_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2279_ _0152_ _0155_ _0160_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__or3_4
XFILLER_0_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1650_ _0819_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__clkbuf_4
X_1581_ _0883_ _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__nor2_2
X_2202_ _1474_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__buf_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2133_ _1402_ _1405_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__or2b_1
X_2064_ top8227.demux.state_machine.currentAddress\[1\] VGND VGND VPWR VPWR _1337_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_71_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2897_ _1407_ _0429_ _0626_ _0703_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__o41a_1
XFILLER_0_44_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1917_ _0823_ _0937_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2966_ _0341_ _0296_ _0763_ _0717_ top8227.internalDataflow.addressLowBusModule.busInputs\[28\]
+ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1779_ _1025_ _1034_ _1041_ _1067_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__or4_1
X_1848_ _1025_ _0978_ _1070_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2820_ _0643_ _0503_ _0644_ _0445_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\]
+ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__a32o_1
X_2751_ _0174_ top8227.internalDataflow.addressLowBusModule.busInputs\[36\] _0593_
+ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2682_ _0135_ _0159_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__nand2_1
X_1633_ _0936_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__nor2_1
X_1564_ _0817_ _0860_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__o21a_1
X_1702_ _1004_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3096_ clknet_4_1_0_clk _0056_ net40 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_2116_ _1378_ _1361_ _1368_ _1373_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__and4b_1
Xfanout37 net44 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
X_2047_ _0923_ _0950_ _0818_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__o21a_1
Xfanout48 net49 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2949_ _0289_ _0291_ _0741_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2803_ gpio[12] _0553_ _0628_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__mux2_1
X_2734_ _0451_ _0313_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2596_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__buf_2
X_1616_ _0850_ _0851_ _0852_ _0853_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__and4_2
X_2665_ _0473_ _0519_ _0521_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__and3_1
X_1547_ _0821_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__buf_2
X_3148_ clknet_4_7_0_clk top8227.pulse_slower.nextEnableState\[1\] net48 VGND VGND
+ VPWR VPWR top8227.pulse_slower.currentEnableState\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3079_ clknet_4_2_0_clk _0039_ net37 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2381_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] _1468_ _1475_
+ _0262_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2450_ _0322_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__inv_2
Xinput5 dataBusIn[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
X_3002_ net78 _0717_ _0789_ _0796_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2717_ _0570_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2648_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] _0457_ VGND
+ VGND VPWR VPWR _0506_ sky130_fd_sc_hd__and2_1
X_2579_ _1399_ _1409_ _0430_ _0437_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1950_ _1088_ _1112_ _1202_ _1215_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1881_ _1119_ _1134_ _1162_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__or3_1
X_2502_ top8227.PSRCurrentValue\[2\] _0368_ _0380_ _0381_ VGND VGND VPWR VPWR _0382_
+ sky130_fd_sc_hd__a31o_1
X_2364_ _1493_ _0245_ _0237_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__o21ai_1
X_2433_ _1305_ _0314_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2295_ _1484_ _1492_ _0176_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2080_ _1348_ _1350_ _1351_ _1352_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__or4b_1
XFILLER_0_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1933_ _0883_ _0834_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__nor2_2
X_2982_ _0351_ _0337_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__nand2_1
X_1864_ _0911_ _0839_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1795_ _0971_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2347_ _1384_ _0225_ _0227_ _0228_ net21 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2416_ _0155_ _0160_ _0152_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__o21a_1
X_2278_ _0139_ _0159_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1580_ _0853_ _0852_ _0851_ _0850_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_53_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2132_ _0929_ _0939_ _1403_ _1404_ _0957_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__a32o_1
X_2201_ _1469_ _1472_ _1467_ _1473_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__and4b_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2063_ _1014_ _0868_ _1335_ _0981_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2896_ _0704_ _0614_ _0705_ _0440_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__or4b_1
XFILLER_0_44_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1847_ _1126_ _1128_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2965_ _0295_ _0288_ _0292_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__nand3_1
X_1916_ _1038_ _1051_ _1056_ _1080_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1778_ _1021_ _1047_ _1056_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2681_ _0201_ _0468_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2750_ _0597_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1701_ _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1632_ _0928_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__clkbuf_4
X_1563_ _0867_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__clkbuf_4
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3095_ clknet_4_0_0_clk _0055_ net35 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_2115_ _1387_ _1381_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__and2_2
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout49 net50 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_4
X_2046_ _1146_ _1151_ _0891_ _1318_ _0955_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__o41a_1
XFILLER_0_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout38 net39 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2879_ _0694_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2948_ _0747_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2802_ _0632_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
X_2664_ _0459_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__nand2_1
X_2733_ _0459_ _0578_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2595_ _0442_ _0426_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__or2_1
X_1546_ top8227.demux.state_machine.currentInstruction\[0\] VGND VGND VPWR VPWR _0851_
+ sky130_fd_sc_hd__clkbuf_4
X_1615_ _0919_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__buf_4
X_3147_ clknet_4_7_0_clk top8227.pulse_slower.nextEnableState\[0\] net43 VGND VGND
+ VPWR VPWR top8227.pulse_slower.currentEnableState\[0\] sky130_fd_sc_hd__dfrtp_1
X_3078_ clknet_4_8_0_clk _0038_ net38 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2029_ top8227.demux.state_machine.currentAddress\[12\] top8227.demux.state_machine.currentAddress\[10\]
+ top8227.demux.state_machine.currentAddress\[4\] _1301_ VGND VGND VPWR VPWR _1302_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2380_ net2 net94 _1469_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
+ _0261_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__a221o_1
Xinput6 dataBusIn[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_4
X_3001_ _0341_ _0792_ _0795_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2647_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] _0459_ VGND
+ VGND VPWR VPWR _0505_ sky130_fd_sc_hd__nor2_1
X_2716_ _0569_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] _0444_
+ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2578_ _1413_ _0434_ _0435_ _0436_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__or4_1
X_1529_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _1145_ _1157_ _1160_ _1161_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2501_ _1247_ _0363_ _0379_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__and3_1
X_2432_ _0310_ _0313_ _1333_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__mux2_2
X_2363_ _1384_ _0225_ _0227_ net21 VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a31oi_4
X_2294_ _0166_ _0173_ _1493_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap24 _0119_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
XFILLER_0_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1932_ _1052_ _1108_ _1169_ _1210_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2981_ _0141_ _0721_ _0775_ _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__a22o_1
X_1863_ _1142_ _1143_ _1144_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__or3_1
X_1794_ _1077_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2415_ _0161_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2277_ _0158_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__buf_2
X_2346_ _1307_ _1333_ _1342_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2131_ _0871_ _0925_ _0920_ _0928_ _1267_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__a311o_1
X_2062_ top8227.branchBackward top8227.branchForward VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__or2_2
X_2200_ _0975_ _1465_ _1458_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__or3_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2964_ _0758_ _0761_ _0341_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2895_ _1016_ _1317_ _1275_ _0987_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__a22o_1
X_1915_ _0823_ _0911_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__nor2_2
X_1846_ _1127_ _1031_ _1062_ _1108_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1777_ top8227.demux.state_machine.currentAddress\[5\] _1035_ _1064_ _1066_ VGND
+ VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2329_ top8227.internalDataflow.accRegToDB\[2\] _1386_ _0210_ VGND VGND VPWR VPWR
+ _0211_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1631_ _0850_ _0853_ _0852_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__or3b_2
XFILLER_0_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2680_ _0191_ _0447_ _0448_ _0190_ _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__a221o_2
XFILLER_0_38_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1700_ _1002_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__buf_2
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1562_ _0861_ _0862_ _0863_ _0866_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__or4b_1
XFILLER_0_39_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2045_ _0941_ _0949_ _1291_ _1317_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__o31a_1
X_3094_ clknet_4_0_0_clk _0054_ net34 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_2114_ _1373_ _1368_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__nand2_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout39 net44 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_4
X_2947_ _0746_ top8227.internalDataflow.addressLowBusModule.busInputs\[26\] _0717_
+ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2878_ _0215_ top8227.internalDataflow.accRegToDB\[2\] net22 VGND VGND VPWR VPWR
+ _0694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1829_ _1040_ _1050_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__and2b_2
XFILLER_0_40_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2801_ gpio[11] _0536_ _0628_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2663_ _0453_ _0511_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__or2_1
X_2732_ _0472_ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__xnor2_1
X_1614_ top8227.demux.state_machine.currentInstruction\[0\] _0821_ _0820_ _0828_ VGND
+ VGND VPWR VPWR _0919_ sky130_fd_sc_hd__or4b_1
X_2594_ _0446_ _0447_ _0448_ _0245_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__a221o_2
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1545_ _0828_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__buf_2
XFILLER_0_22_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3077_ clknet_4_6_0_clk _0037_ net42 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_1
X_3146_ clknet_4_2_0_clk _0106_ net34 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_2028_ top8227.demux.state_machine.currentAddress\[3\] top8227.demux.state_machine.currentAddress\[11\]
+ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__or2_2
XFILLER_0_9_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput7 dataBusIn[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_4
X_3000_ _0323_ _0794_ _0731_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2646_ net75 _0445_ _0475_ _0477_ _0504_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__a221o_1
X_2715_ _0561_ _0562_ _0567_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2577_ _0971_ _1419_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1528_ top8227.demux.state_machine.currentInstruction\[1\] top8227.demux.state_machine.currentInstruction\[0\]
+ top8227.demux.state_machine.currentInstruction\[2\] top8227.demux.state_machine.currentInstruction\[3\]
+ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__or4b_1
XFILLER_0_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3129_ clknet_4_1_0_clk _0089_ net40 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2431_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _1468_ _1475_
+ _0312_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2500_ _1247_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__nand2_1
X_2293_ _1305_ _0174_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__nand2_1
X_2362_ _0243_ _0139_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2629_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] _0455_ VGND VGND
+ VPWR VPWR _0488_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2980_ _0355_ _0315_ _0301_ _0730_ _0731_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__o221a_1
XFILLER_0_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1931_ _1209_ _1033_ _1055_ _1085_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__a22o_1
X_1793_ top8227.demux.state_machine.currentAddress\[9\] _1076_ _0979_ VGND VGND VPWR
+ VPWR _1077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1862_ _0872_ _1033_ _1098_ net26 VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__a22o_1
X_2414_ _0288_ _0292_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2276_ _0127_ _0157_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__or2_1
X_2345_ top8227.internalDataflow.accRegToDB\[0\] _1386_ _1388_ top8227.internalDataflow.stackBusModule.busInputs\[40\]
+ _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2130_ _0936_ _0928_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__or2_1
X_2061_ _1285_ _1306_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1914_ _1038_ _1057_ _1085_ _1033_ _0890_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2963_ _0182_ _0721_ _0759_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1845_ _0912_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__buf_4
X_2894_ _1447_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1776_ _1034_ _1065_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2328_ top8227.internalDataflow.stackBusModule.busInputs\[34\] _1380_ _1388_ top8227.internalDataflow.stackBusModule.busInputs\[42\]
+ _0209_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2259_ _1483_ _0140_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1630_ _0931_ _0932_ _0933_ _0934_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1561_ _0864_ _0834_ _0846_ _0865_ _0825_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__a41o_1
XFILLER_0_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2044_ _1316_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__clkbuf_4
X_2113_ _1385_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__clkbuf_4
X_3093_ clknet_4_3_0_clk _0053_ net35 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_2877_ _0693_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
X_2946_ _0740_ _0745_ _0341_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1828_ _0937_ _0885_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__nor2_1
X_1759_ net5 _1017_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__nand2_2
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2731_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\] _0582_ VGND
+ VGND VPWR VPWR _0583_ sky130_fd_sc_hd__xor2_1
X_2800_ _0631_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1544_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__clkbuf_4
X_2662_ _0453_ _0465_ _0511_ _0458_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__a31o_1
X_1613_ _0888_ _0900_ _0910_ _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__or4_2
X_2593_ _0449_ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3145_ clknet_4_2_0_clk _0105_ net34 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2027_ _1285_ _1293_ _1299_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__or3_1
X_3076_ clknet_4_2_0_clk _0036_ net34 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2929_ _1246_ _1296_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__nand2_2
XFILLER_0_32_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 dataBusIn[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_0_19_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2714_ _0564_ _0566_ _0425_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2645_ _0501_ _0502_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__and3_1
X_2576_ top8227.demux.state_machine.timeState\[1\] _0916_ _0912_ _0915_ VGND VGND
+ VPWR VPWR _0435_ sky130_fd_sc_hd__o22a_1
X_1527_ top8227.demux.state_machine.currentInstruction\[5\] VGND VGND VPWR VPWR _0832_
+ sky130_fd_sc_hd__clkbuf_4
X_3128_ clknet_4_1_0_clk _0088_ net40 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3059_ clknet_4_12_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
+ net39 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2430_ net8 net25 _1469_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\]
+ _0311_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__a221o_1
X_2361_ _0240_ _0242_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__nor2_2
X_2292_ _0168_ _0173_ _1333_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__mux2_2
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2559_ _0419_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
X_2628_ _0485_ _0455_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap26 _1102_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
XFILLER_0_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1930_ _0911_ _0834_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__nor2_4
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1792_ _1060_ _1064_ _1065_ _1075_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__a31o_1
X_1861_ _0891_ _1092_ _1055_ _1098_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__a22o_1
X_2344_ top8227.internalDataflow.stackBusModule.busInputs\[32\] _1380_ _1391_ top8227.internalDataflow.addressLowBusModule.busInputs\[24\]
+ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a22o_1
X_2413_ _0182_ _0294_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__nand2_1
X_2275_ top8227.internalDataflow.addressLowBusModule.busInputs\[29\] _0130_ _0132_
+ net6 _0156_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_59_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ _1332_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__clkbuf_4
X_2893_ _0436_ _0700_ _0701_ _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1913_ _0855_ _0979_ _1053_ _1085_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__a2bb2o_1
X_2962_ _0355_ _0152_ _0293_ _0730_ _0731_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1844_ _0905_ _1031_ _1072_ _1108_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__a22o_1
X_1775_ _1041_ _1050_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2327_ top8227.internalDataflow.addressLowBusModule.busInputs\[34\] _1390_ _1391_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[26\] VGND VGND VPWR VPWR
+ _0209_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2258_ _1495_ _0135_ _0139_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2189_ _1461_ _1444_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1560_ _0828_ top8227.demux.state_machine.currentInstruction\[0\] _0821_ _0820_ VGND
+ VGND VPWR VPWR _0865_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_55_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2112_ _1378_ _1361_ _1368_ _1373_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__and4bb_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2043_ _0907_ top8227.demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR _1316_
+ sky130_fd_sc_hd__or2_1
X_3092_ clknet_4_0_0_clk _0052_ net35 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2876_ _0271_ top8227.internalDataflow.accRegToDB\[1\] _0691_ VGND VGND VPWR VPWR
+ _0693_ sky130_fd_sc_hd__mux2_1
X_1827_ _0886_ _1032_ _1057_ _1108_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a22o_1
X_2945_ _0289_ _0744_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1689_ _0990_ _0991_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1758_ net2 _1048_ _1050_ _1035_ net58 VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2730_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\] _0459_ _0581_
+ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2661_ _0213_ _0447_ _0448_ _0212_ _0517_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__a221o_2
XFILLER_0_41_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1543_ _0832_ _0835_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__nor2_1
X_1612_ _0912_ _0914_ _0915_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__o31a_1
X_2592_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3075_ clknet_4_8_0_clk _0035_ net38 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
X_3144_ clknet_4_2_0_clk _0104_ net37 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2026_ _1252_ _1297_ _1298_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__or3_1
X_2859_ _0484_ _0498_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2928_ _0282_ _0280_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 nrst VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_2713_ _0564_ _0566_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__or2_1
X_2644_ _0476_ _0443_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__nor2_4
XFILLER_0_42_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2575_ _0914_ _0431_ _0432_ _0896_ _0433_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a221o_1
X_1526_ _0827_ _0830_ _0826_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__or3_1
X_3127_ clknet_4_1_0_clk _0087_ net40 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3058_ clknet_4_12_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
+ net39 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[0\] sky130_fd_sc_hd__dfrtp_4
X_2009_ _1003_ _1281_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2291_ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] _1468_ _1475_
+ _0172_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a211o_1
X_2360_ top8227.internalDataflow.addressLowBusModule.busInputs\[24\] _0130_ _0132_
+ net1 _0241_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2627_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] _0456_ VGND VGND
+ VPWR VPWR _0486_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2558_ net16 _1494_ _0412_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
X_1509_ top8227.demux.state_machine.timeState\[2\] VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__clkbuf_4
X_2489_ _0943_ _0944_ _0952_ _1005_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__o31a_1
XFILLER_0_69_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap27 net28 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1860_ _1135_ _1092_ _1038_ _1141_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1791_ _1020_ _1073_ _1074_ _1072_ net2 VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__a32o_1
X_2343_ top8227.internalDataflow.addressLowBusModule.busInputs\[32\] _1390_ VGND VGND
+ VPWR VPWR _0225_ sky130_fd_sc_hd__nand2_1
X_2274_ top8227.internalDataflow.addressLowBusModule.busInputs\[37\] net24 _0125_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] _0126_ VGND VGND VPWR
+ VPWR _0156_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2412_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1989_ _0907_ _0957_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2892_ _1005_ _1009_ _0916_ _1400_ _1127_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__o41a_1
XFILLER_0_56_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1912_ _1192_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
X_1843_ _0862_ _1034_ _1053_ _1103_ _1124_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__a221o_1
X_2961_ _0295_ _0722_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__or2_1
X_1774_ _1025_ _1047_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2326_ _1331_ _0207_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2257_ _0138_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2188_ _0890_ _1250_ _1001_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 top8227.instructionLoader.interruptInjector.irqSync.nextQ2 VGND VGND VPWR VPWR
+ net51 sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ clknet_4_6_0_clk _0051_ net43 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_2111_ _1383_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__buf_4
X_3160_ clknet_4_2_0_clk VGND VGND VPWR VPWR gpio[23] sky130_fd_sc_hd__buf_2
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2042_ _1175_ _1090_ _1314_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2875_ _0692_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2944_ _0726_ _0742_ _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1826_ _0978_ _1019_ _1107_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__and3_2
X_1688_ _0814_ _0859_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__and2b_1
X_1757_ net7 _1049_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__nor2_1
X_2309_ net4 _1434_ _1435_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\]
+ net19 VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1611_ top8227.demux.state_machine.timeState\[5\] VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2660_ _0207_ _0451_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2591_ _1312_ _0447_ _1493_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__or3b_1
X_1542_ _0826_ _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3074_ clknet_4_7_0_clk _0034_ net48 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
X_2025_ _1003_ _0868_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__and2_2
X_3143_ clknet_4_2_0_clk _0103_ net37 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2927_ _1261_ _0726_ _0290_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2858_ _0675_ _0677_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__nand2_1
X_2789_ _1212_ _0887_ _1400_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1809_ _1030_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__clkbuf_4
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2643_ _0480_ _0500_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__nand2_1
X_2574_ _0818_ _0898_ _0951_ _1316_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__a22o_1
X_2712_ _0146_ _0447_ _0448_ _0145_ _0565_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1525_ _0829_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__clkbuf_4
X_3057_ clknet_4_14_0_clk _0025_ net49 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2008_ _0839_ _0846_ _0879_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__a21oi_1
X_3126_ clknet_4_3_0_clk _0086_ net39 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2290_ top8227.internalDataflow.accRegToDB\[4\] _1478_ _1469_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\]
+ _0171_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2626_ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] VGND VGND VPWR
+ VPWR _0485_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2557_ _0418_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2488_ _1295_ _1325_ _1015_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3109_ clknet_4_1_0_clk _0069_ net40 VGND VGND VPWR VPWR gpio[10] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1790_ _1060_ _1056_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2411_ _0175_ _0181_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__and2_1
X_2342_ _0216_ _0223_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__xnor2_4
X_2273_ _0139_ _0154_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1988_ _1259_ _1260_ top8227.PSRCurrentValue\[3\] VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__or3b_4
X_2609_ _0466_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__nor2_1
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2960_ _0295_ _0288_ _0757_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2891_ _1009_ _1273_ _0432_ _1096_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__o31a_1
XFILLER_0_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1842_ _0849_ _0856_ _1032_ _1024_ _1053_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__a32o_1
X_1911_ _1119_ _1191_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__or2_1
X_1773_ _1055_ _1057_ _1059_ _1063_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2187_ _1271_ _1443_ _1459_ _0972_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__o31a_1
X_2325_ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] _1468_ _1475_
+ _0206_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__a211oi_1
X_2256_ _1245_ _0137_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2110_ _1380_ _1381_ _1382_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__or3_1
X_3090_ clknet_4_1_0_clk _0050_ net35 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[32\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold2 top8227.instructionLoader.interruptInjector.nmiSync.nextQ2 VGND VGND VPWR VPWR
+ net52 sky130_fd_sc_hd__dlygate4sd3_1
X_2041_ _0908_ _0994_ _0997_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2943_ _0290_ _0741_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__and2_1
X_2874_ _0238_ top8227.internalDataflow.accRegToDB\[0\] _0691_ VGND VGND VPWR VPWR
+ _0692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1756_ _1021_ _1017_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__nand2_2
X_1825_ _1021_ net7 _1018_ _1040_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__and4bb_2
X_1687_ _0907_ _0818_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__nor2_1
X_2308_ _0188_ _0189_ _0165_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2239_ gpio[19] _0981_ top8227.pulse_slower.nextEnableState\[0\] _0120_ VGND VGND
+ VPWR VPWR _0121_ sky130_fd_sc_hd__and4_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1610_ _0874_ _0846_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__nor2_2
X_2590_ _0235_ _0236_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1541_ _0845_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__buf_2
X_3142_ clknet_4_2_0_clk _0102_ net39 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2024_ _0955_ _1294_ _1295_ _1003_ _1296_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__a221o_1
X_3073_ clknet_4_8_0_clk net52 net38 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2857_ _0471_ _0676_ _0459_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__o21ai_1
X_2926_ _1261_ _0290_ _0726_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2788_ _1013_ _0618_ _0619_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__a211o_1
X_1808_ _0871_ _0928_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1739_ _1033_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__clkbuf_4
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2711_ _0451_ _0150_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2642_ _0480_ _0500_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__or2_1
X_2573_ top8227.demux.state_machine.timeState\[5\] top8227.demux.state_machine.timeState\[3\]
+ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__or2_1
X_1524_ _0828_ _0820_ _0821_ top8227.demux.state_machine.currentInstruction\[0\] VGND
+ VGND VPWR VPWR _0829_ sky130_fd_sc_hd__or4bb_1
X_3125_ clknet_4_1_0_clk _0085_ net40 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3056_ clknet_4_14_0_clk _0024_ net49 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2007_ _1278_ _1279_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2909_ _0135_ _0712_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2625_ _0482_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2487_ _1247_ _0359_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__nand2_1
X_2556_ net86 _0153_ _0412_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3108_ clknet_4_5_0_clk _0068_ net41 VGND VGND VPWR VPWR gpio[9] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3039_ clknet_4_10_0_clk _0011_ net47 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2341_ _0218_ _0222_ _0139_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__mux2_2
X_2410_ _0204_ _0286_ _0289_ _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__o22ai_2
X_2272_ _1484_ _1492_ _0153_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1987_ _1078_ _0985_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2608_ _0279_ _0243_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__nand2_1
X_2539_ top8227.PSRCurrentValue\[2\] top8227.demux.setInterruptFlag top8227.instructionLoader.interruptInjector.irqGenerated
+ top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ VGND
+ VGND VPWR VPWR _0407_ sky130_fd_sc_hd__or4b_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2890_ _1014_ _0620_ _1321_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1910_ _1145_ _1171_ _1183_ _1190_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__or4_1
XFILLER_0_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1841_ _1120_ _1092_ _1080_ net26 _1122_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1772_ _1038_ _1060_ _1062_ _1034_ net91 VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__a32o_1
X_2324_ net3 net25 _1469_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\]
+ _0205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__a221o_1
X_2186_ _0896_ _0912_ _1002_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__o21a_1
X_2255_ _0955_ _1321_ _0136_ _1298_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2040_ top8227.demux.state_machine.currentAddress\[12\] _1262_ _0971_ VGND VGND VPWR
+ VPWR _1313_ sky130_fd_sc_hd__a21oi_1
Xhold3 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning VGND
+ VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2873_ _0372_ _0689_ _0690_ _1247_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__o31ai_4
X_2942_ _0290_ _0741_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1824_ _0849_ _0921_ _1032_ _1101_ _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__a311o_1
X_1686_ top8227.demux.state_machine.currentAddress\[6\] _0988_ VGND VGND VPWR VPWR
+ _0989_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1755_ _0977_ _1047_ _1025_ _0986_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2238_ top8227.demux.state_machine.currentAddress\[5\] _0987_ _1001_ VGND VGND VPWR
+ VPWR _0120_ sky130_fd_sc_hd__o21a_1
X_2307_ top8227.internalDataflow.accRegToDB\[3\] _1386_ _1384_ VGND VGND VPWR VPWR
+ _0189_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2169_ _1343_ _1396_ _1441_ _1342_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1540_ top8227.demux.state_machine.currentInstruction\[0\] top8227.demux.state_machine.currentInstruction\[2\]
+ top8227.demux.state_machine.currentInstruction\[3\] top8227.demux.state_machine.currentInstruction\[1\]
+ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3141_ clknet_4_2_0_clk _0101_ net37 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_2023_ _1003_ _0891_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__and2_2
X_3072_ clknet_4_2_0_clk top8227.instructionLoader.interruptInjector.nmiSync.in net37
+ VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiSync.nextQ2 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2856_ _0157_ _0470_ _0135_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__a21oi_1
X_1807_ _1081_ _1083_ _1088_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2925_ _0204_ _0286_ _0292_ _0287_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2787_ top8227.demux.state_machine.timeState\[3\] _1096_ _1127_ _0620_ _0982_ VGND
+ VGND VPWR VPWR _0621_ sky130_fd_sc_hd__a221o_1
X_1669_ _0869_ _0918_ _0956_ _0972_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1738_ _1032_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2710_ _0554_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2641_ _0481_ _0484_ _0498_ _0482_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__a311o_1
X_2572_ _0859_ top8227.demux.state_machine.timeState\[1\] top8227.demux.state_machine.timeState\[5\]
+ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__or3_1
X_1523_ top8227.demux.state_machine.currentInstruction\[1\] VGND VGND VPWR VPWR _0828_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3055_ clknet_4_15_0_clk _0023_ net49 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3124_ clknet_4_3_0_clk _0084_ net39 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2006_ _1003_ _0894_ _0901_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2908_ gpio[6] _0708_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__nand2_1
X_2839_ _0427_ _0469_ _0180_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2624_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] _0456_ VGND VGND
+ VPWR VPWR _0483_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2486_ _1247_ _1257_ _0357_ _0367_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2555_ _0417_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap19 _1440_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
X_3107_ clknet_4_1_0_clk _0067_ net40 VGND VGND VPWR VPWR gpio[8] sky130_fd_sc_hd__dfrtp_4
X_3038_ clknet_4_11_0_clk _0010_ net45 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2271_ _0145_ _0150_ _1493_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__mux2_2
X_2340_ top8227.demux.nmi _0219_ _0221_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_55_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1986_ _1248_ _1258_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2607_ _0222_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2469_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__inv_2
X_2538_ top8227.demux.nmi _0405_ _0406_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1840_ _1020_ _1103_ _1113_ _1091_ _1121_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1771_ _1061_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__clkbuf_4
X_2323_ top8227.internalDataflow.accRegToDB\[2\] _1478_ _1476_ top8227.PSRCurrentValue\[2\]
+ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__a22o_1
X_2254_ _1004_ _1127_ _1184_ _1014_ _1288_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2185_ _0981_ _1445_ _1451_ _1457_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__o22a_2
X_1969_ _1244_ VGND VGND VPWR VPWR top8227.pulse_slower.nextEnableState\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 top8227.demux.state_machine.currentAddress\[8\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2872_ _0931_ _0952_ _1006_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2941_ _1484_ _1259_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__nor2_2
X_1823_ _1037_ _1072_ _1080_ _1104_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__a31o_1
X_1754_ net4 _1043_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__or2_2
XFILLER_0_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1685_ _0987_ top8227.demux.state_machine.currentAddress\[12\] VGND VGND VPWR VPWR
+ _0988_ sky130_fd_sc_hd__nor2_1
X_2237_ _1497_ _1506_ _0118_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__nor3_1
X_2306_ top8227.internalDataflow.stackBusModule.busInputs\[35\] _1380_ _1388_ top8227.internalDataflow.stackBusModule.busInputs\[43\]
+ _0187_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a221o_1
X_2168_ net7 _1434_ _1435_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\]
+ net19 VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2099_ _0981_ _1369_ _1371_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3071_ clknet_4_15_0_clk net51 net50 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3140_ clknet_4_8_0_clk _0100_ net38 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_2022_ _0871_ _0876_ _0920_ _0825_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_10_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2786_ _1015_ _0431_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2855_ _0135_ _0463_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__a21o_1
X_1806_ _0894_ _1084_ _1031_ _1085_ _1087_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2924_ net74 _0717_ _0720_ _0725_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__a22o_1
X_1599_ _0903_ _0897_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__and2_2
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1668_ gpio[19] _0968_ top8227.pulse_slower.nextEnableState\[0\] _0971_ VGND VGND
+ VPWR VPWR _0972_ sky130_fd_sc_hd__o211a_4
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1737_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__buf_2
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2640_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _0456_ VGND VGND
+ VPWR VPWR _0499_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2571_ _1013_ _0816_ _0428_ _1274_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o41a_1
X_1522_ top8227.PSRCurrentValue\[0\] VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2005_ top8227.demux.state_machine.timeState\[1\] _0849_ _0894_ VGND VGND VPWR VPWR
+ _1278_ sky130_fd_sc_hd__and3_1
X_3054_ clknet_4_14_0_clk _0022_ net49 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3123_ clknet_4_3_0_clk _0083_ net36 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_2907_ _0159_ _0711_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2838_ _0458_ _0462_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2769_ net72 _0193_ _0605_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__mux2_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2623_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] _0456_ VGND VGND
+ VPWR VPWR _0482_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2554_ net14 _0176_ _0412_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__mux2_1
X_2485_ _0358_ _0361_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3106_ clknet_4_8_0_clk _0066_ net45 VGND VGND VPWR VPWR top8227.demux.reset sky130_fd_sc_hd__dfrtp_4
X_3037_ clknet_4_14_0_clk _0009_ net46 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2270_ _1305_ _0151_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1985_ _0907_ _1158_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2606_ _0320_ _0464_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2537_ top8227.demux.nmi top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning
+ top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI VGND
+ VGND VPWR VPWR _0406_ sky130_fd_sc_hd__or3b_1
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2399_ _0272_ _0280_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__xnor2_4
X_2468_ _0342_ net30 net23 _1491_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__a31o_2
XFILLER_0_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1770_ _1042_ _1043_ _1051_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2253_ _0127_ _0134_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__or2_2
X_2184_ _1453_ _1374_ _1456_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__nor3_1
X_2322_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1968_ top8227.pulse_slower.currentEnableState\[1\] net64 VGND VGND VPWR VPWR _1244_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1899_ _0883_ _0920_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 top8227.instructionLoader.interruptInjector.resetDetected VGND VGND VPWR VPWR
+ net55 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2940_ _0350_ _0289_ _0739_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__o21ba_1
X_2871_ _1209_ _0942_ _0951_ _1015_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__o31a_1
XFILLER_0_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1753_ net60 _1035_ _1046_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a21o_1
X_1822_ _0944_ _1030_ _1102_ _1103_ _1059_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__a221o_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1684_ top8227.demux.state_machine.currentAddress\[1\] VGND VGND VPWR VPWR _0987_
+ sky130_fd_sc_hd__clkbuf_4
X_2167_ _1434_ _1435_ _1438_ _1439_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__nor4_1
X_2236_ net27 _1508_ _0975_ _1424_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__a211oi_2
X_2305_ top8227.internalDataflow.addressLowBusModule.busInputs\[35\] _1390_ _1391_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[27\] VGND VGND VPWR VPWR
+ _0187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2098_ _1175_ _1314_ _1370_ _0993_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3070_ clknet_4_15_0_clk top8227.instructionLoader.interruptInjector.interruptRequest
+ net50 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.irqSync.nextQ2
+ sky130_fd_sc_hd__dfrtp_1
X_2021_ _0883_ _0936_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__nor2_2
XFILLER_0_57_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2923_ _0259_ _0721_ _0723_ _0724_ _0351_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_72_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2785_ _1005_ _1009_ _0916_ _1184_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__o32a_1
X_2854_ _0472_ _0464_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1805_ _1057_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__and2_2
X_1736_ _1030_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__clkbuf_4
X_1598_ _0835_ _0832_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__and2b_2
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1667_ top8227.demux.isAddressing net33 VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__nand2_4
XFILLER_0_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _1485_ _1489_ _1491_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__a21o_2
XFILLER_0_48_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2570_ _0868_ _1273_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3122_ clknet_4_7_0_clk _0082_ net43 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_1521_ _0825_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3053_ clknet_4_15_0_clk _0021_ net49 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2004_ _1184_ _1273_ _1276_ _0982_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__a211o_1
X_2906_ gpio[5] _0708_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1719_ _1013_ _1010_ _1012_ _1014_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a22o_1
X_2699_ _0541_ _0542_ _0536_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__mux2_1
X_2837_ _0201_ _0461_ _0180_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__o21a_1
X_2768_ _0608_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2622_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _0456_ VGND VGND
+ VPWR VPWR _0481_ sky130_fd_sc_hd__or2_1
X_2553_ _0416_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2484_ _0362_ _0363_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__mux2_1
X_3105_ clknet_4_3_0_clk _0065_ net34 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_3036_ clknet_4_10_0_clk _0008_ net46 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_73_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1984_ _1252_ _1253_ _1255_ _1256_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2605_ _0134_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__or2_1
X_2467_ _1005_ _0949_ _1251_ _1256_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2536_ net67 _0404_ _0405_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2398_ _0275_ _0279_ _0139_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__mux2_2
XFILLER_0_46_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3019_ _0806_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2321_ _0195_ _0202_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2183_ _0859_ _0915_ _1309_ _1454_ _1455_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__a2111o_1
X_2252_ top8227.internalDataflow.addressLowBusModule.busInputs\[30\] _0130_ _0132_
+ net7 _0133_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1967_ _1243_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
X_1898_ _0826_ _0920_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2519_ _0395_ VGND VGND VPWR VPWR gpio[24] sky130_fd_sc_hd__buf_1
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 top8227.branchForward VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
X_2870_ _0688_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1683_ _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__buf_4
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1752_ _1025_ _0979_ _1045_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__and3_1
X_1821_ _1040_ _1050_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__and2_2
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _1331_ _0185_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2166_ _1013_ _1009_ _1096_ _1245_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__o211ai_2
X_2235_ _1419_ _1507_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__and2_1
X_2097_ top8227.demux.state_machine.currentAddress\[11\] top8227.demux.state_machine.currentAddress\[12\]
+ top8227.demux.state_machine.currentAddress\[4\] _0971_ VGND VGND VPWR VPWR _1370_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2999_ _0324_ _0793_ _0722_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2020_ _1253_ _1286_ _1290_ _1292_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__or4_1
X_2853_ _0673_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2922_ _1247_ _1296_ _0249_ _0272_ _0354_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__a32o_1
X_2784_ _0835_ _0894_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1666_ top8227.demux.state_machine.currentAddress\[8\] top8227.demux.state_machine.currentAddress\[0\]
+ top8227.demux.state_machine.currentAddress\[2\] top8227.demux.state_machine.currentAddress\[9\]
+ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__nor4_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1804_ net29 _1041_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__nor2_2
X_1735_ _0976_ _0977_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__or2_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ _0894_ _0901_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__and2_2
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2149_ _1001_ _1263_ _0971_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__a21oi_2
X_2218_ _1447_ _1450_ _1490_ _0976_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1520_ _0824_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3121_ clknet_4_5_0_clk _0081_ net42 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3052_ clknet_4_15_0_clk _0020_ net49 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_2003_ _0914_ _1275_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__and2_1
X_2905_ _0180_ _0710_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__nand2_1
X_2836_ _0658_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1718_ _0916_ _1010_ _1012_ _1009_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2698_ _0167_ _0447_ _0448_ _0166_ _0552_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__a221o_2
X_1649_ _0941_ _0945_ _0948_ _0953_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__or4_1
X_2767_ net68 _0215_ _0605_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__mux2_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2621_ _0478_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__nor2_1
X_2552_ net13 _0196_ _0412_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2483_ _0898_ _0905_ _0364_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3104_ clknet_4_0_0_clk _0064_ net35 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_3035_ clknet_4_10_0_clk _0007_ net45 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2819_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _0642_ VGND VGND
+ VPWR VPWR _0644_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2604_ _0159_ _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__or2b_1
X_1983_ _0872_ _1158_ _1005_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2466_ _1357_ _0346_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2535_ _0380_ _0363_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__nand2b_1
X_2397_ _0219_ _0276_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__o21ba_2
X_3018_ top8227.internalDataflow.stackBusModule.busInputs\[38\] _1482_ _0799_ VGND
+ VGND VPWR VPWR _0806_ sky130_fd_sc_hd__mux2_1
Xwire31 _0343_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2251_ top8227.internalDataflow.addressLowBusModule.busInputs\[38\] net24 _0125_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] _0126_ VGND VGND VPWR
+ VPWR _0133_ sky130_fd_sc_hd__a221o_1
X_2320_ _0197_ _0201_ _0139_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
X_2182_ _0815_ _1321_ _1278_ _0981_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__a211o_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1966_ _1238_ _1240_ _1242_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1897_ _0923_ _1092_ _1054_ _1080_ _1177_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__a221o_1
X_2518_ clknet_4_6_0_clk top8227.pulse_slower.nextEnableState\[0\] VGND VGND VPWR
+ VPWR _0395_ sky130_fd_sc_hd__and2_2
XFILLER_0_59_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2449_ _0325_ _0326_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold7 top8227.branchBackward VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
X_1820_ _0976_ net29 _1041_ _1073_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__nor4_2
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1682_ _0984_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1751_ _1041_ _1044_ _1026_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__o21ai_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _0860_ _1274_ _0868_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__o21ai_1
X_2303_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] _1468_ _1475_
+ _0184_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2165_ _1322_ _1436_ _1437_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__or3_1
X_2096_ _1110_ _1135_ _0948_ _1214_ _0993_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__o41a_1
XFILLER_0_63_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1949_ _1226_ _1033_ _1055_ _1111_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2998_ _0322_ _0730_ _0258_ _0354_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_31_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2852_ _0672_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] _0444_
+ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2783_ _1508_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__inv_2
X_1803_ _1040_ _1023_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__and2b_2
X_2921_ _0718_ _0722_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__nor2_1
X_1665_ _0969_ VGND VGND VPWR VPWR top8227.pulse_slower.nextEnableState\[0\] sky130_fd_sc_hd__inv_2
X_1596_ _0832_ _0835_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__and2b_2
X_1734_ _1029_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2217_ top8227.demux.state_machine.currentAddress\[12\] _1275_ VGND VGND VPWR VPWR
+ _1490_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2079_ _0859_ _0896_ _0914_ _0814_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__a22oi_1
X_2148_ _0817_ _1420_ _0868_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3120_ clknet_4_4_0_clk _0080_ net42 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_3051_ clknet_4_6_0_clk _0026_ net43 VGND VGND VPWR VPWR top8227.branchForward sky130_fd_sc_hd__dfrtp_1
X_2002_ _0819_ _1274_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__or2_2
X_2904_ gpio[4] _0708_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__nand2_1
X_2835_ _0657_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] _0444_
+ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2766_ _0607_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1717_ _1015_ _1010_ _1012_ _1006_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__a22o_1
X_1579_ _0883_ _0842_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__nor2_4
X_2697_ _0451_ _0173_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__and2b_1
X_1648_ _0949_ _0950_ _0951_ _0952_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__or4_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2620_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] _0456_ VGND
+ VGND VPWR VPWR _0479_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2551_ _0415_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
X_2482_ _1267_ _1260_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__nor2_4
X_3103_ clknet_4_0_0_clk _0063_ net35 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_3034_ clknet_4_11_0_clk _0006_ net45 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2818_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _0642_ VGND VGND
+ VPWR VPWR _0643_ sky130_fd_sc_hd__nand2_1
X_2749_ _0193_ top8227.internalDataflow.addressLowBusModule.busInputs\[35\] _0593_
+ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__mux2_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1982_ _1254_ _0923_ _1004_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2603_ _0179_ _0201_ _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__nor3_1
XFILLER_0_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2534_ _1010_ _1018_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__nor2_1
X_2396_ top8227.internalDataflow.addressLowBusModule.busInputs\[25\] _0130_ _0132_
+ net2 _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__a221o_1
X_2465_ _1005_ _0923_ _1282_ _0982_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3017_ _0805_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2250_ _0131_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2181_ _0815_ _0886_ _0950_ _0993_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1965_ _1185_ _1194_ _1228_ _1241_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2517_ _0394_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
+ sky130_fd_sc_hd__clkbuf_1
X_1896_ _1175_ _1176_ _0978_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__mux2_1
X_2379_ top8227.internalDataflow.accRegToDB\[1\] _1478_ _1476_ top8227.PSRCurrentValue\[1\]
+ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__a22o_1
X_2448_ _0304_ _0327_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_61_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold8 top8227.demux.state_machine.currentAddress\[3\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1750_ _1042_ _1043_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1681_ _0969_ _0983_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2164_ _1294_ _0896_ _1002_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__o21a_1
X_2302_ net4 net25 _1469_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\]
+ _0183_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__a221o_1
X_2233_ _0985_ _1501_ _1505_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2095_ _0969_ _0983_ _1367_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__or3_2
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1948_ _0937_ _0925_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1879_ _1020_ _1103_ _1130_ _1033_ _0924_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2997_ _0338_ _0790_ _0791_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2920_ _1209_ _0364_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__nand2_4
X_2851_ _0667_ _0671_ _0425_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1802_ _0832_ _0835_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__and2_1
X_2782_ _1263_ _1265_ _1273_ _0615_ _1078_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__a221o_1
X_1733_ _1016_ _1028_ _0979_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__mux2_1
X_1664_ top8227.pulse_slower.currentEnableState\[1\] top8227.pulse_slower.currentEnableState\[0\]
+ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__or2_2
X_1595_ _0815_ _0889_ _0892_ _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__a211o_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2147_ _1001_ _0955_ _0859_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__or3_1
X_2216_ _1335_ _1270_ _1486_ _1004_ _1488_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2078_ _1151_ _0902_ top8227.demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR
+ _1351_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3050_ clknet_4_13_0_clk _0019_ net49 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_2001_ _0908_ _0815_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__or2_2
X_2903_ _0201_ _0709_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1716_ net73 _1010_ _1012_ _0916_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__a22o_1
X_2834_ _0653_ _0654_ _0656_ _0477_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__a22o_1
X_2696_ _0531_ _0549_ _0548_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__o21ai_1
X_2765_ top8227.internalDataflow.stackBusModule.busInputs\[41\] _0271_ _0605_ VGND
+ VGND VPWR VPWR _0607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1647_ _0901_ _0897_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__and2_2
X_1578_ _0874_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__buf_4
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2550_ net79 _0217_ _0412_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2481_ _0916_ top8227.demux.setInterruptFlag _1078_ _1096_ _0832_ VGND VGND VPWR
+ VPWR _0363_ sky130_fd_sc_hd__a41o_1
XFILLER_0_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3102_ clknet_4_0_0_clk _0062_ net34 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_3033_ clknet_4_10_0_clk _0005_ net47 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2817_ _0491_ _0490_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__and2b_1
X_2679_ _0185_ _0451_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__nor2_1
X_2748_ _0596_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1981_ _1195_ _1135_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2533_ net82 _0986_ _0389_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__o21ba_1
X_2602_ _0222_ _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2395_ top8227.internalDataflow.addressLowBusModule.busInputs\[33\] net24 _0125_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] VGND VGND VPWR VPWR
+ _0277_ sky130_fd_sc_hd__a22o_1
X_2464_ _1279_ _0344_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or3_1
X_3016_ net92 _0151_ _0799_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__mux2_1
Xwire33 _0970_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
XFILLER_0_73_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2180_ _0868_ _1308_ _1452_ _1001_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1964_ _1109_ _1126_ _1165_ _1168_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1895_ _1040_ _1018_ _1027_ _1047_ _1069_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_59_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2447_ _0300_ _0328_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__nand2_2
X_2516_ _0390_ _0391_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or3b_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2378_ _0249_ _0258_ _0259_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__a21o_2
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 top8227.demux.state_machine.currentAddress\[0\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1680_ _0971_ _0968_ gpio[19] VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__a21oi_2
X_2301_ top8227.internalDataflow.accRegToDB\[3\] _1478_ _1476_ top8227.PSRCurrentValue\[3\]
+ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2232_ _1270_ _1503_ _1504_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__or3_1
X_2163_ _1127_ _0887_ _0955_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2094_ _1362_ _1363_ _1366_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1947_ _1221_ _1222_ _1223_ _1224_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__or4_1
X_1878_ _1158_ _1034_ _1024_ _1055_ _1159_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2996_ _0338_ _0790_ _0350_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2850_ _0668_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__xnor2_1
X_1663_ _0964_ _0930_ _0966_ _0967_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__o31a_2
X_2781_ _1016_ _1317_ _1266_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1801_ _0914_ _1031_ _1062_ _1082_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1732_ _1020_ _1024_ _1027_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__a21oi_1
X_1594_ top8227.demux.state_machine.timeState\[3\] _0896_ _0898_ _0819_ VGND VGND
+ VPWR VPWR _0899_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2077_ _0814_ _0890_ _0891_ top8227.demux.state_machine.timeState\[4\] _1349_ VGND
+ VGND VPWR VPWR _1350_ sky130_fd_sc_hd__a221o_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2146_ _0950_ _1317_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__nand2_1
X_2215_ _0914_ _1274_ _1280_ _1487_ _1251_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_63_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2979_ _0303_ _0722_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2000_ _0960_ _0990_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__nand2_2
XFILLER_0_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2902_ gpio[3] _0708_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__nand2_1
X_2833_ _0201_ _0655_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1715_ _1014_ _1010_ _1012_ _1015_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a22o_1
X_2695_ _0531_ _0548_ _0549_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__or3_1
X_1646_ _0883_ _0865_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__nor2_2
X_2764_ _0606_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1577_ _0872_ _0877_ _0880_ _0881_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__or4_2
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2129_ _1400_ _0880_ _0941_ _1316_ _1401_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__a221o_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2480_ _1246_ _1257_ _0361_ _0827_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_23_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3101_ clknet_4_3_0_clk _0061_ net36 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_3032_ clknet_4_12_0_clk _0004_ net45 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2816_ _0639_ _0640_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2678_ _0530_ _0531_ _0532_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__or3b_1
X_1629_ _0928_ _0865_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__nor2_2
XFILLER_0_41_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2747_ _0215_ top8227.internalDataflow.addressLowBusModule.busInputs\[34\] _0593_
+ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1980_ _0877_ _1212_ _1151_ _1003_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__o31a_1
X_2601_ _0279_ _0243_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__or2_1
X_2463_ _1005_ _1009_ _0965_ _1096_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__o31a_1
X_2532_ top8227.demux.nmi _0381_ _0403_ net53 VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2394_ top8227.demux.nmi top8227.demux.reset VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__and2b_1
X_3015_ _0804_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire23 _0349_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1894_ _0937_ _0920_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__nor2_1
X_1963_ _1133_ _1239_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2446_ _0299_ _0182_ _0296_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__nand3_1
X_2515_ _0338_ _0392_ _0339_ top8227.PSRCurrentValue\[3\] _0386_ VGND VGND VPWR VPWR
+ _0393_ sky130_fd_sc_hd__a2111o_1
X_2377_ _0244_ _0248_ _0239_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _1498_ _1321_ _1347_ _0981_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2300_ _0175_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__or2_2
X_2162_ _0985_ _1432_ _1425_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2093_ _1364_ _1365_ top8227.demux.state_machine.currentAddress\[3\] _0971_ VGND
+ VGND VPWR VPWR _1366_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2995_ _0324_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1946_ _1170_ _1178_ _1189_ _1203_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__or4_1
X_1877_ _0877_ _1031_ _1085_ _1102_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__a22o_1
X_2429_ top8227.internalDataflow.accRegToDB\[7\] _1478_ _1476_ top8227.PSRCurrentValue\[7\]
+ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1800_ _0978_ _1019_ _1024_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__and3_1
X_1662_ _0907_ _0929_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__or2_1
X_2780_ _1006_ top8227.demux.state_machine.currentAddress\[5\] _1301_ _1262_ _1499_
+ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1731_ _1025_ _1026_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__or2_1
X_1593_ _0849_ _0897_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__and2_2
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _1013_ _1184_ _1289_ _0982_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2076_ top8227.demux.state_machine.timeState\[4\] top8227.demux.state_machine.timeState\[6\]
+ top8227.demux.state_machine.timeState\[1\] _0901_ _0856_ VGND VGND VPWR VPWR _1349_
+ sky130_fd_sc_hd__o311a_1
X_2145_ _1399_ _1409_ _1413_ _1417_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__nor4_1
XFILLER_0_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1929_ _1089_ _1106_ _1129_ _1157_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2978_ net69 _0717_ _0770_ _0774_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2832_ _0466_ _0467_ _0539_ _0461_ _0458_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__o32a_1
XFILLER_0_42_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2763_ top8227.internalDataflow.stackBusModule.busInputs\[40\] _0238_ _0605_ VGND
+ VGND VPWR VPWR _0606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2901_ gpio[2] _0708_ _0466_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__a21o_1
X_2694_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] _0457_ _0532_
+ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__o21a_1
X_1576_ _0839_ _0834_ _0874_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__a21oi_2
X_1645_ _0825_ _0885_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__nor2_4
X_1714_ _0955_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__clkbuf_4
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2128_ _0846_ _0842_ _0885_ _0911_ _0957_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__a311oi_1
X_2059_ _1312_ _1331_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__and2b_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3100_ clknet_4_3_0_clk _0060_ net35 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_3031_ clknet_4_10_0_clk _0000_ net47 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2815_ _0467_ _0460_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__nand2_1
X_2746_ _0595_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2677_ _0530_ _0531_ _0532_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__o21bai_1
X_1628_ _0852_ _0853_ _0832_ _0835_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__and4b_1
X_1559_ _0828_ _0851_ _0821_ _0820_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_41_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2600_ _0458_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2462_ _1184_ _1273_ _1420_ _1127_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__a22o_1
X_2531_ top8227.demux.nmi _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__or2_1
X_2393_ _1484_ _1492_ _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3014_ net87 _0174_ _0799_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2729_ _0571_ _0572_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1962_ _1101_ _1122_ _1201_ _1227_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1893_ _0847_ _0979_ _1053_ _1098_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__a2bb2o_1
X_2376_ _1271_ _0255_ _0257_ _0985_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__o211a_1
X_2445_ _0303_ _0161_ _0300_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__nand3_1
X_2514_ _0323_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _1014_ _0912_ _1184_ _1009_ _1502_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__a221o_1
X_2161_ _1433_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__buf_2
XFILLER_0_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2092_ top8227.demux.state_machine.currentAddress\[5\] _1090_ top8227.demux.state_machine.currentAddress\[10\]
+ _1267_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__a211o_1
X_1945_ _1095_ _1104_ _1123_ _1210_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2994_ _0341_ _0788_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1876_ _0826_ _0876_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2428_ _1343_ _0308_ _0309_ _1342_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a22o_1
X_2359_ top8227.internalDataflow.addressLowBusModule.busInputs\[32\] net24 _0125_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] VGND VGND VPWR VPWR
+ _0241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1592_ _0851_ _0852_ _0853_ _0850_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__and4b_1
X_1661_ _0872_ _0877_ _0880_ _0881_ _0965_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__o41a_1
XFILLER_0_40_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1730_ net4 net3 _1018_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__nand3_1
X_2144_ _0981_ _0899_ _1414_ _1416_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__or4_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _1184_ _0950_ _1291_ _1411_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__or4_1
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2075_ _0814_ _0889_ _0915_ top8227.demux.state_machine.timeState\[6\] _1347_ VGND
+ VGND VPWR VPWR _1348_ sky130_fd_sc_hd__a221o_1
X_1928_ _1207_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2977_ _1261_ _0772_ _0773_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__or3_1
X_1859_ net7 _1049_ _1062_ _1138_ _1140_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__o311a_1
XFILLER_0_12_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2900_ gpio[1] _0708_ _0279_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__a21bo_1
X_2831_ _0493_ _0646_ _0652_ _0425_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__o31a_1
X_1713_ _0815_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2762_ _0604_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2693_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] _0457_ VGND
+ VGND VPWR VPWR _0548_ sky130_fd_sc_hd__xor2_1
X_1575_ _0830_ _0839_ _0879_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__a21oi_1
X_1644_ _0879_ _0885_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__nor2_4
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ _0814_ _0859_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__or2_2
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2058_ _1313_ _1315_ _1330_ _0976_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__a211o_4
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3030_ _0813_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2676_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] _0457_ _0527_
+ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__a21o_1
X_2814_ _0243_ _0472_ _0539_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2745_ _0271_ top8227.internalDataflow.addressLowBusModule.busInputs\[33\] _0593_
+ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1627_ _0928_ _0842_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__nor2_2
X_1558_ _0839_ _0842_ _0825_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__a21oi_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3159_ clknet_4_12_0_clk _0117_ net44 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2530_ top8227.PSRCurrentValue\[2\] top8227.demux.setInterruptFlag _1010_ VGND VGND
+ VPWR VPWR _0402_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2392_ _1331_ _0263_ _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__a21oi_2
X_2461_ _1005_ _1411_ _1276_ _1292_ _1248_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire25 net94 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
X_3013_ _0803_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2659_ net90 _0445_ _0509_ _0503_ _0516_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2728_ net76 _0445_ _0573_ _0503_ _0580_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1892_ _1172_ _1092_ _1053_ _1164_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1961_ _1083_ _1095_ _1232_ _1237_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__or4_1
XFILLER_0_70_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2513_ _0387_ _1494_ _1247_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__and3b_1
X_2375_ _1004_ _0987_ top8227.freeCarry _0256_ _1355_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2444_ _0141_ _0304_ _0324_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _0985_ _1425_ _1432_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap1 _1395_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_1
X_2091_ _0907_ top8227.demux.state_machine.currentAddress\[1\] _1016_ top8227.demux.state_machine.currentAddress\[11\]
+ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1944_ _1081_ _1128_ _1132_ _1150_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2993_ _0330_ _0771_ _0787_ _0784_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__a31o_1
X_1875_ _1150_ _1155_ _1156_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2427_ _1021_ _1434_ _1435_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\]
+ net19 VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
X_2289_ net5 _1477_ _1476_ _0170_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2358_ _1013_ _1245_ _1278_ _0126_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__and4b_1
XFILLER_0_66_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1591_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__clkbuf_4
X_1660_ top8227.demux.state_machine.timeState\[4\] _0814_ VGND VGND VPWR VPWR _0965_
+ sky130_fd_sc_hd__or2_2
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2143_ top8227.demux.state_machine.timeState\[5\] _0915_ _0951_ _1317_ _1415_ VGND
+ VGND VPWR VPWR _1416_ sky130_fd_sc_hd__a221o_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _1004_ _0884_ _1287_ _1297_ _1282_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2074_ _0850_ top8227.demux.state_machine.timeState\[4\] _0903_ _1346_ VGND VGND
+ VPWR VPWR _1347_ sky130_fd_sc_hd__and4_1
X_1927_ _1118_ _1134_ _1206_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__or3_1
X_2976_ _0329_ _0331_ _0771_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__and3_1
X_1858_ _1139_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__inv_2
X_1789_ _1070_ _1062_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__or2_2
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2830_ _0493_ _0646_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2692_ _0547_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
X_1712_ _1009_ _1010_ _1012_ _1013_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 _0704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1643_ _0946_ _0947_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__or2_1
X_2761_ _1246_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1574_ _0878_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__buf_4
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ _0960_ _1397_ _1317_ _1398_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__a2bb2o_1
X_2057_ _1319_ _1329_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__nor2_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2959_ _0351_ _0335_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__nand2_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2813_ _0443_ _0638_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2675_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] _0457_ VGND
+ VGND VPWR VPWR _0531_ sky130_fd_sc_hd__and2_1
X_1626_ _0864_ _0885_ _0928_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2744_ _0594_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1557_ _0830_ _0825_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__nor2_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ clknet_4_4_0_clk _0049_ net41 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2109_ _1373_ _1361_ _1368_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__and3_1
X_3158_ clknet_4_10_0_clk _0116_ net46 VGND VGND VPWR VPWR top8227.demux.isAddressing
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_17_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2460_ _1270_ _1298_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2391_ _1331_ _0268_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3012_ net70 _0193_ _0799_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2658_ _0425_ _0515_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__nor2_1
X_1609_ _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__clkbuf_4
X_2727_ _0425_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__nor2_1
X_2589_ _0447_ _1312_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1891_ _0826_ _0842_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1960_ _1181_ _1198_ _1235_ _1236_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2512_ top8227.PSRCurrentValue\[6\] _0386_ _0388_ _0389_ top8227.negEdgeDetector.q1
+ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2443_ _0141_ _0304_ _0324_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a21oi_1
X_2374_ _1337_ _0996_ _1263_ _1262_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2090_ _0908_ top8227.demux.state_machine.currentAddress\[1\] _1090_ _1317_ _0980_
+ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__o311a_1
Xmax_cap2 _1477_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2992_ _0781_ _0329_ _0741_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__or3b_1
XFILLER_0_61_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1874_ _1037_ _1052_ _1080_ _1031_ _0840_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__a32o_1
X_1943_ _1114_ _1142_ _1161_ _1167_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__or4_1
X_2426_ _1384_ _0307_ net20 VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2288_ _1014_ _1096_ _0169_ _1294_ _1003_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2357_ _1305_ _0238_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1590_ _0848_ _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__and2_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2142_ _0859_ top8227.demux.state_machine.timeState\[5\] _0912_ VGND VGND VPWR VPWR
+ _1415_ sky130_fd_sc_hd__o21a_1
X_2073_ _0853_ _0852_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__and2b_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _1248_ _1255_ _1245_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2975_ _0331_ _0771_ _0329_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__a21oi_1
X_1926_ _1171_ _1200_ _1204_ _1205_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1788_ net77 _1035_ _1055_ _1072_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__a22o_1
X_1857_ _1080_ _1103_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__or2_1
X_2409_ _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2691_ _0546_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] _0444_
+ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__mux2_1
X_1711_ _0859_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_2 top8227.PSRCurrentValue\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
X_1642_ _0879_ _0846_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__nor2_1
X_2760_ _1015_ _0948_ _0602_ _1006_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1573_ _0832_ _0835_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__or2b_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ _0819_ _0927_ _0945_ _0891_ _0923_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__a2111o_1
X_2056_ _1323_ _1324_ _1326_ _1328_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__or4_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1909_ _1185_ _1189_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__or2_1
X_2958_ top8227.internalDataflow.addressLowBusModule.busInputs\[27\] _0717_ _0750_
+ _0752_ _0756_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2889_ _0699_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2812_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _0637_ _0477_
+ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__mux2_1
X_2743_ _0238_ top8227.internalDataflow.addressLowBusModule.busInputs\[32\] _0593_
+ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2674_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] _0458_ VGND
+ VGND VPWR VPWR _0530_ sky130_fd_sc_hd__nor2_1
X_1625_ _0929_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__inv_2
X_1556_ _0823_ _0825_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3157_ clknet_4_6_0_clk _0115_ net43 VGND VGND VPWR VPWR top8227.branchBackward sky130_fd_sc_hd__dfrtp_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3088_ clknet_4_4_0_clk _0048_ net41 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[22\]
+ sky130_fd_sc_hd__dfrtp_2
X_2039_ _1298_ _1311_ _0972_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__o21ai_4
X_2108_ _1373_ _1378_ _1361_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3011_ _0802_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
X_2390_ _1305_ _0271_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__and2_2
XFILLER_0_58_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2726_ _0576_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2657_ _0511_ _0514_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__xnor2_1
X_1608_ _0903_ _0894_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__and2_1
X_2588_ _1245_ _1334_ _1340_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__a21o_2
X_1539_ top8227.PSRCurrentValue\[1\] _0840_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1890_ _1166_ _1168_ _1170_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__or3_1
X_2511_ gpio[20] _1010_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__nor2_2
XFILLER_0_59_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2373_ _1324_ _0252_ _0253_ _0254_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2442_ _0322_ _0323_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2709_ _0458_ _0553_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1942_ _1220_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2991_ net63 _0717_ _0780_ _0786_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1873_ _1154_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__inv_2
X_2356_ _1333_ _0229_ _0233_ _0237_ _1312_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__o32a_2
X_2425_ top8227.internalDataflow.accRegToDB\[7\] _1386_ _0306_ VGND VGND VPWR VPWR
+ _0307_ sky130_fd_sc_hd__a21oi_1
X_2287_ top8227.demux.reset top8227.demux.nmi top8227.demux.setInterruptFlag VGND
+ VGND VPWR VPWR _0169_ sky130_fd_sc_hd__nor3_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _1305_ _1482_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2141_ top8227.demux.state_machine.timeState\[1\] top8227.demux.state_machine.timeState\[5\]
+ _0914_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__o21a_1
X_2072_ _1320_ _1344_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__or2_1
X_1925_ _0861_ _1034_ _1053_ _1111_ _1173_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2974_ _0332_ _0333_ _0323_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1787_ _1071_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__clkbuf_4
X_1856_ _1060_ _1062_ _1137_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2339_ top8227.internalDataflow.addressLowBusModule.busInputs\[26\] _0130_ _0132_
+ net3 _0220_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a221o_1
X_2408_ _0260_ _0281_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2690_ _0425_ _0533_ _0534_ _0545_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__a31o_1
X_1710_ _1011_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__clkbuf_2
X_1572_ _0874_ _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__nor2_2
XANTENNA_3 top8227.PSRCurrentValue\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1641_ _0911_ _0842_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2124_ _0872_ _0877_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__nor2_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2055_ _0934_ _1295_ _1327_ _0818_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__o31a_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2888_ _0314_ top8227.internalDataflow.accRegToDB\[7\] net22 VGND VGND VPWR VPWR
+ _0699_ sky130_fd_sc_hd__mux2_1
X_1839_ _0830_ _0937_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1908_ _1187_ _1188_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__or2_1
X_2957_ _0287_ _0731_ _0755_ _0350_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2811_ _0243_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__inv_2
X_2742_ _1247_ _0592_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__nand2_4
XFILLER_0_26_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2673_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] _0445_ _0523_
+ _0477_ _0529_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__a221o_1
X_1624_ _0871_ _0925_ _0920_ _0928_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__a31o_1
X_1555_ _0819_ _0837_ _0844_ _0858_ _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__a41o_1
X_3087_ clknet_4_4_0_clk _0047_ net41 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[21\]
+ sky130_fd_sc_hd__dfrtp_2
X_2107_ _1379_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__clkbuf_4
X_3156_ clknet_4_2_0_clk _0114_ net34 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2038_ _1002_ _1308_ _1309_ _1310_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3010_ net83 _0215_ _0799_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire28 _1418_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
XFILLER_0_73_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2656_ _0459_ _0512_ _0513_ _0473_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__o211a_1
X_2725_ _1441_ _0447_ _0448_ _1396_ _0577_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__a221o_2
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2587_ _0231_ _0232_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__or2_1
X_1607_ _0911_ _0864_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__nor2_4
X_1538_ _0826_ _0842_ top8227.PSRCurrentValue\[1\] VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3139_ clknet_4_9_0_clk _0099_ net39 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2510_ _0924_ _0364_ _0387_ _1260_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2372_ _0982_ _1255_ _1282_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2441_ _0315_ _0321_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__nor2_2
X_2639_ _0485_ _0472_ _0486_ _0496_ _0497_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__o221ai_4
X_2708_ _0557_ _0558_ _0560_ _0476_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1941_ _1166_ _1190_ _1204_ _1219_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2990_ _0331_ _0771_ _0783_ _0785_ _1261_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__a311oi_1
X_1872_ _1151_ _1030_ _1153_ _0977_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2286_ _1343_ _0166_ _0167_ _1342_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__a22o_1
X_2355_ _0235_ _0236_ _1331_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__nand3b_2
X_2424_ top8227.internalDataflow.stackBusModule.busInputs\[39\] _1380_ _1388_ top8227.internalDataflow.stackBusModule.busInputs\[47\]
+ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2140_ _0819_ _0906_ _1410_ _1412_ _0909_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__a2111o_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2071_ _0941_ _0949_ _1291_ _1281_ _0818_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__o41a_1
X_1924_ _1201_ _1202_ _1203_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2973_ _0351_ _0336_ _0766_ _0769_ _0341_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__a311o_1
X_1855_ _1064_ _1097_ _1136_ _1036_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1786_ _1025_ _1070_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__and2_1
X_2269_ _0147_ _0150_ _1333_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__mux2_2
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2338_ top8227.internalDataflow.addressLowBusModule.busInputs\[34\] net24 _0125_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] VGND VGND VPWR VPWR
+ _0220_ sky130_fd_sc_hd__a22o_1
X_2407_ _0224_ _0284_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__xor2_4
XFILLER_0_62_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold40 top8227.internalDataflow.addressHighBusModule.busInputs\[17\] VGND VGND VPWR
+ VPWR net90 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1571_ _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__clkbuf_4
X_1640_ _0942_ _0943_ _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2123_ _1384_ _1394_ net20 VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__a21oi_2
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2054_ _0850_ _0851_ _0933_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1838_ _0830_ _0911_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2887_ _0698_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
X_1907_ _1020_ _1113_ _1164_ _1032_ _0947_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2956_ _0203_ _0722_ _0754_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__o21ai_1
X_1769_ _1049_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2672_ _0527_ _0503_ _0528_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__and3b_1
X_2810_ _0636_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
X_2741_ _1348_ _1496_ _0591_ _1352_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__or4b_2
XFILLER_0_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1554_ top8227.demux.state_machine.timeState\[6\] VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__buf_2
X_1623_ _0832_ _0835_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__nand2_4
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

