VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO silly_synthesizer
  CLASS BLOCK ;
  FOREIGN silly_synthesizer ;
  ORIGIN 0.000 0.000 ;
  SIZE 228.665 BY 239.385 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 224.665 217.640 228.665 218.240 ;
    END
  END cs
  PIN gpio[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 235.385 206.450 239.385 ;
    END
  END gpio[0]
  PIN gpio[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 235.385 119.510 239.385 ;
    END
  END gpio[10]
  PIN gpio[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END gpio[11]
  PIN gpio[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END gpio[12]
  PIN gpio[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.665 34.040 228.665 34.640 ;
    END
  END gpio[13]
  PIN gpio[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END gpio[14]
  PIN gpio[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.665 170.040 228.665 170.640 ;
    END
  END gpio[15]
  PIN gpio[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END gpio[16]
  PIN gpio[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gpio[1]
  PIN gpio[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END gpio[2]
  PIN gpio[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END gpio[3]
  PIN gpio[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 235.385 74.430 239.385 ;
    END
  END gpio[4]
  PIN gpio[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.665 125.840 228.665 126.440 ;
    END
  END gpio[5]
  PIN gpio[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END gpio[6]
  PIN gpio[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 161.090 235.385 161.370 239.385 ;
    END
  END gpio[7]
  PIN gpio[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END gpio[8]
  PIN gpio[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END gpio[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 235.385 32.570 239.385 ;
    END
  END nrst
  PIN pwm
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.665 78.240 228.665 78.840 ;
    END
  END pwm
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 228.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 228.720 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 223.100 228.565 ;
      LAYER met1 ;
        RECT 0.070 10.640 223.490 228.720 ;
      LAYER met2 ;
        RECT 0.100 235.105 32.010 235.385 ;
        RECT 32.850 235.105 73.870 235.385 ;
        RECT 74.710 235.105 118.950 235.385 ;
        RECT 119.790 235.105 160.810 235.385 ;
        RECT 161.650 235.105 205.890 235.385 ;
        RECT 206.730 235.105 223.470 235.385 ;
        RECT 0.100 4.280 223.470 235.105 ;
        RECT 0.650 3.670 41.670 4.280 ;
        RECT 42.510 3.670 86.750 4.280 ;
        RECT 87.590 3.670 128.610 4.280 ;
        RECT 129.450 3.670 173.690 4.280 ;
        RECT 174.530 3.670 215.550 4.280 ;
        RECT 216.390 3.670 223.470 4.280 ;
      LAYER met3 ;
        RECT 4.400 227.440 224.665 228.645 ;
        RECT 4.000 218.640 224.665 227.440 ;
        RECT 4.000 217.240 224.265 218.640 ;
        RECT 4.000 184.640 224.665 217.240 ;
        RECT 4.400 183.240 224.665 184.640 ;
        RECT 4.000 171.040 224.665 183.240 ;
        RECT 4.000 169.640 224.265 171.040 ;
        RECT 4.000 137.040 224.665 169.640 ;
        RECT 4.400 135.640 224.665 137.040 ;
        RECT 4.000 126.840 224.665 135.640 ;
        RECT 4.000 125.440 224.265 126.840 ;
        RECT 4.000 92.840 224.665 125.440 ;
        RECT 4.400 91.440 224.665 92.840 ;
        RECT 4.000 79.240 224.665 91.440 ;
        RECT 4.000 77.840 224.265 79.240 ;
        RECT 4.000 45.240 224.665 77.840 ;
        RECT 4.400 43.840 224.665 45.240 ;
        RECT 4.000 35.040 224.665 43.840 ;
        RECT 4.000 33.640 224.265 35.040 ;
        RECT 4.000 10.715 224.665 33.640 ;
      LAYER met4 ;
        RECT 52.735 26.695 97.440 154.185 ;
        RECT 99.840 26.695 156.105 154.185 ;
  END
END silly_synthesizer
END LIBRARY

