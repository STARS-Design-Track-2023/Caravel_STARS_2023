magic
tech sky130A
magscale 1 2
timestamp 1691529709
<< obsli1 >>
rect 1104 2159 41400 42449
<< obsm1 >>
rect 14 2128 41938 42560
<< metal2 >>
rect 3238 43864 3294 44664
rect 7102 43864 7158 44664
rect 10966 43864 11022 44664
rect 14830 43864 14886 44664
rect 18694 43864 18750 44664
rect 22558 43864 22614 44664
rect 26422 43864 26478 44664
rect 30286 43864 30342 44664
rect 34150 43864 34206 44664
rect 38014 43864 38070 44664
rect 41878 43864 41934 44664
rect 18 0 74 800
rect 3882 0 3938 800
rect 7746 0 7802 800
rect 11610 0 11666 800
rect 15474 0 15530 800
rect 19338 0 19394 800
rect 23202 0 23258 800
rect 27066 0 27122 800
rect 30930 0 30986 800
rect 34794 0 34850 800
rect 38658 0 38714 800
<< obsm2 >>
rect 20 43808 3182 44305
rect 3350 43808 7046 44305
rect 7214 43808 10910 44305
rect 11078 43808 14774 44305
rect 14942 43808 18638 44305
rect 18806 43808 22502 44305
rect 22670 43808 26366 44305
rect 26534 43808 30230 44305
rect 30398 43808 34094 44305
rect 34262 43808 37958 44305
rect 38126 43808 41822 44305
rect 20 856 41932 43808
rect 130 31 3826 856
rect 3994 31 7690 856
rect 7858 31 11554 856
rect 11722 31 15418 856
rect 15586 31 19282 856
rect 19450 31 23146 856
rect 23314 31 27010 856
rect 27178 31 30874 856
rect 31042 31 34738 856
rect 34906 31 38602 856
rect 38770 31 41932 856
<< metal3 >>
rect 0 44208 800 44328
rect 41720 40808 42520 40928
rect 0 40128 800 40248
rect 41720 36728 42520 36848
rect 0 36048 800 36168
rect 41720 32648 42520 32768
rect 0 31968 800 32088
rect 41720 28568 42520 28688
rect 0 27888 800 28008
rect 41720 24488 42520 24608
rect 0 23808 800 23928
rect 41720 20408 42520 20528
rect 0 19728 800 19848
rect 41720 16328 42520 16448
rect 0 15648 800 15768
rect 41720 12248 42520 12368
rect 0 11568 800 11688
rect 41720 8168 42520 8288
rect 0 7488 800 7608
rect 41720 4088 42520 4208
rect 0 3408 800 3528
rect 41720 8 42520 128
<< obsm3 >>
rect 880 44128 41720 44301
rect 800 41008 41720 44128
rect 800 40728 41640 41008
rect 800 40328 41720 40728
rect 880 40048 41720 40328
rect 800 36928 41720 40048
rect 800 36648 41640 36928
rect 800 36248 41720 36648
rect 880 35968 41720 36248
rect 800 32848 41720 35968
rect 800 32568 41640 32848
rect 800 32168 41720 32568
rect 880 31888 41720 32168
rect 800 28768 41720 31888
rect 800 28488 41640 28768
rect 800 28088 41720 28488
rect 880 27808 41720 28088
rect 800 24688 41720 27808
rect 800 24408 41640 24688
rect 800 24008 41720 24408
rect 880 23728 41720 24008
rect 800 20608 41720 23728
rect 800 20328 41640 20608
rect 800 19928 41720 20328
rect 880 19648 41720 19928
rect 800 16528 41720 19648
rect 800 16248 41640 16528
rect 800 15848 41720 16248
rect 880 15568 41720 15848
rect 800 12448 41720 15568
rect 800 12168 41640 12448
rect 800 11768 41720 12168
rect 880 11488 41720 11768
rect 800 8368 41720 11488
rect 800 8088 41640 8368
rect 800 7688 41720 8088
rect 880 7408 41720 7688
rect 800 4288 41720 7408
rect 800 4008 41640 4288
rect 800 3608 41720 4008
rect 880 3328 41720 3608
rect 800 208 41720 3328
rect 800 35 41640 208
<< metal4 >>
rect 4208 2128 4528 42480
rect 19568 2128 19888 42480
rect 34928 2128 35248 42480
<< obsm4 >>
rect 5027 2619 19488 41853
rect 19968 2619 31221 41853
<< labels >>
rlabel metal3 s 0 15648 800 15768 6 M10ClkOut
port 1 nsew signal output
rlabel metal4 s 19568 2128 19888 42480 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 42480 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 42480 6 VPWR
port 3 nsew power bidirectional
rlabel metal2 s 38658 0 38714 800 6 addressBusHigh[0]
port 4 nsew signal output
rlabel metal2 s 18694 43864 18750 44664 6 addressBusHigh[1]
port 5 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 addressBusHigh[2]
port 6 nsew signal output
rlabel metal3 s 41720 8168 42520 8288 6 addressBusHigh[3]
port 7 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 addressBusHigh[4]
port 8 nsew signal output
rlabel metal3 s 41720 4088 42520 4208 6 addressBusHigh[5]
port 9 nsew signal output
rlabel metal3 s 41720 8 42520 128 6 addressBusHigh[6]
port 10 nsew signal output
rlabel metal3 s 41720 32648 42520 32768 6 addressBusHigh[7]
port 11 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 addressBusLow[0]
port 12 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 addressBusLow[1]
port 13 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 addressBusLow[2]
port 14 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 addressBusLow[3]
port 15 nsew signal output
rlabel metal3 s 41720 36728 42520 36848 6 addressBusLow[4]
port 16 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 addressBusLow[5]
port 17 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 addressBusLow[6]
port 18 nsew signal output
rlabel metal2 s 38014 43864 38070 44664 6 addressBusLow[7]
port 19 nsew signal output
rlabel metal2 s 26422 43864 26478 44664 6 clk
port 20 nsew signal input
rlabel metal3 s 41720 24488 42520 24608 6 dataBusEnable
port 21 nsew signal input
rlabel metal2 s 34150 43864 34206 44664 6 dataBusInput[0]
port 22 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 dataBusInput[1]
port 23 nsew signal input
rlabel metal3 s 41720 40808 42520 40928 6 dataBusInput[2]
port 24 nsew signal input
rlabel metal2 s 7102 43864 7158 44664 6 dataBusInput[3]
port 25 nsew signal input
rlabel metal2 s 18 0 74 800 6 dataBusInput[4]
port 26 nsew signal input
rlabel metal2 s 22558 43864 22614 44664 6 dataBusInput[5]
port 27 nsew signal input
rlabel metal3 s 41720 28568 42520 28688 6 dataBusInput[6]
port 28 nsew signal input
rlabel metal2 s 3238 43864 3294 44664 6 dataBusInput[7]
port 29 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 dataBusOutput[0]
port 30 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 dataBusOutput[1]
port 31 nsew signal output
rlabel metal2 s 30286 43864 30342 44664 6 dataBusOutput[2]
port 32 nsew signal output
rlabel metal3 s 41720 12248 42520 12368 6 dataBusOutput[3]
port 33 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 dataBusOutput[4]
port 34 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 dataBusOutput[5]
port 35 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 dataBusOutput[6]
port 36 nsew signal output
rlabel metal3 s 41720 16328 42520 16448 6 dataBusOutput[7]
port 37 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 dataBusSelect
port 38 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 functionalClockOut
port 39 nsew signal output
rlabel metal2 s 41878 43864 41934 44664 6 interruptRequest
port 40 nsew signal input
rlabel metal2 s 10966 43864 11022 44664 6 nonMaskableInterrupt
port 41 nsew signal input
rlabel metal2 s 14830 43864 14886 44664 6 nrst
port 42 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 readNotWrite
port 43 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 ready
port 44 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 setOverflow
port 45 nsew signal input
rlabel metal3 s 41720 20408 42520 20528 6 sync
port 46 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 42520 44664
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6240152
string GDS_FILE /home/designer-25/CUP/openlane/outel8227/runs/23_08_08_14_15/results/signoff/top8227.magic.gds
string GDS_START 1134918
<< end >>

